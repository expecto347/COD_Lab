
`timescale 1ns / 1ps
module cache_tb();

localparam INDEX_WIDTH          = 3;
localparam WORD_OFFSET_WIDTH    = 4;
localparam TOTAL_WORD_NUM       = 1024;

// cache test
reg [31:0]  i_addr_rom [TOTAL_WORD_NUM];
reg [31:0]  d_addr_rom [TOTAL_WORD_NUM];
reg [31:0]  data_ram [TOTAL_WORD_NUM];
reg         wvalid_rom [TOTAL_WORD_NUM];
reg [31:0]  wdata_rom [TOTAL_WORD_NUM];
reg [31:0]  i_test_index = 0;
reg [31:0]  d_test_index = 0;
reg clk = 1'b1, rstn = 1'b0;

initial #5 rstn = 1'b1; 
always #1 clk = ~clk;

// generate data_ram
initial begin
    data_ram[    0] = 'h00000000; 	    data_ram[    1] = 'h00000001; 	    data_ram[    2] = 'h00000002; 	    data_ram[    3] = 'h00000003; 	    data_ram[    4] = 'h00000004; 	    data_ram[    5] = 'h00000005; 	    data_ram[    6] = 'h00000006; 	    data_ram[    7] = 'h00000007; 	
    data_ram[    8] = 'h00000008; 	    data_ram[    9] = 'h00000009; 	    data_ram[   10] = 'h0000000a; 	    data_ram[   11] = 'h0000000b; 	    data_ram[   12] = 'h0000000c; 	    data_ram[   13] = 'h0000000d; 	    data_ram[   14] = 'h0000000e; 	    data_ram[   15] = 'h0000000f; 	
    data_ram[   16] = 'h00000010; 	    data_ram[   17] = 'h00000011; 	    data_ram[   18] = 'h00000012; 	    data_ram[   19] = 'h00000013; 	    data_ram[   20] = 'h00000014; 	    data_ram[   21] = 'h00000015; 	    data_ram[   22] = 'h00000016; 	    data_ram[   23] = 'h00000017; 	
    data_ram[   24] = 'h00000018; 	    data_ram[   25] = 'h00000019; 	    data_ram[   26] = 'h0000001a; 	    data_ram[   27] = 'h0000001b; 	    data_ram[   28] = 'h0000001c; 	    data_ram[   29] = 'h0000001d; 	    data_ram[   30] = 'h0000001e; 	    data_ram[   31] = 'h0000001f; 	
    data_ram[   32] = 'h00000020; 	    data_ram[   33] = 'h00000021; 	    data_ram[   34] = 'h00000022; 	    data_ram[   35] = 'h00000023; 	    data_ram[   36] = 'h00000024; 	    data_ram[   37] = 'h00000025; 	    data_ram[   38] = 'h00000026; 	    data_ram[   39] = 'h00000027; 	
    data_ram[   40] = 'h00000028; 	    data_ram[   41] = 'h00000029; 	    data_ram[   42] = 'h0000002a; 	    data_ram[   43] = 'h0000002b; 	    data_ram[   44] = 'h0000002c; 	    data_ram[   45] = 'h0000002d; 	    data_ram[   46] = 'h0000002e; 	    data_ram[   47] = 'h0000002f; 	
    data_ram[   48] = 'h00000030; 	    data_ram[   49] = 'h00000031; 	    data_ram[   50] = 'h00000032; 	    data_ram[   51] = 'h00000033; 	    data_ram[   52] = 'h00000034; 	    data_ram[   53] = 'h00000035; 	    data_ram[   54] = 'h00000036; 	    data_ram[   55] = 'h00000037; 	
    data_ram[   56] = 'h00000038; 	    data_ram[   57] = 'h00000039; 	    data_ram[   58] = 'h0000003a; 	    data_ram[   59] = 'h0000003b; 	    data_ram[   60] = 'h0000003c; 	    data_ram[   61] = 'h0000003d; 	    data_ram[   62] = 'h0000003e; 	    data_ram[   63] = 'h0000003f; 	
    data_ram[   64] = 'h00000040; 	    data_ram[   65] = 'h00000041; 	    data_ram[   66] = 'h00000042; 	    data_ram[   67] = 'h00000043; 	    data_ram[   68] = 'h00000044; 	    data_ram[   69] = 'h00000045; 	    data_ram[   70] = 'h00000046; 	    data_ram[   71] = 'h00000047; 	
    data_ram[   72] = 'h00000048; 	    data_ram[   73] = 'h00000049; 	    data_ram[   74] = 'h0000004a; 	    data_ram[   75] = 'h0000004b; 	    data_ram[   76] = 'h0000004c; 	    data_ram[   77] = 'h0000004d; 	    data_ram[   78] = 'h0000004e; 	    data_ram[   79] = 'h0000004f; 	
    data_ram[   80] = 'h00000050; 	    data_ram[   81] = 'h00000051; 	    data_ram[   82] = 'h00000052; 	    data_ram[   83] = 'h00000053; 	    data_ram[   84] = 'h00000054; 	    data_ram[   85] = 'h00000055; 	    data_ram[   86] = 'h00000056; 	    data_ram[   87] = 'h00000057; 	
    data_ram[   88] = 'h00000058; 	    data_ram[   89] = 'h00000059; 	    data_ram[   90] = 'h0000005a; 	    data_ram[   91] = 'h0000005b; 	    data_ram[   92] = 'h0000005c; 	    data_ram[   93] = 'h0000005d; 	    data_ram[   94] = 'h0000005e; 	    data_ram[   95] = 'h0000005f; 	
    data_ram[   96] = 'h00000060; 	    data_ram[   97] = 'h00000061; 	    data_ram[   98] = 'h00000062; 	    data_ram[   99] = 'h00000063; 	    data_ram[  100] = 'h00000064; 	    data_ram[  101] = 'h00000065; 	    data_ram[  102] = 'h00000066; 	    data_ram[  103] = 'h00000067; 	
    data_ram[  104] = 'h00000068; 	    data_ram[  105] = 'h00000069; 	    data_ram[  106] = 'h0000006a; 	    data_ram[  107] = 'h0000006b; 	    data_ram[  108] = 'h0000006c; 	    data_ram[  109] = 'h0000006d; 	    data_ram[  110] = 'h0000006e; 	    data_ram[  111] = 'h0000006f; 	
    data_ram[  112] = 'h00000070; 	    data_ram[  113] = 'h00000071; 	    data_ram[  114] = 'h00000072; 	    data_ram[  115] = 'h00000073; 	    data_ram[  116] = 'h00000074; 	    data_ram[  117] = 'h00000075; 	    data_ram[  118] = 'h00000076; 	    data_ram[  119] = 'h00000077; 	
    data_ram[  120] = 'h00000078; 	    data_ram[  121] = 'h00000079; 	    data_ram[  122] = 'h0000007a; 	    data_ram[  123] = 'h0000007b; 	    data_ram[  124] = 'h0000007c; 	    data_ram[  125] = 'h0000007d; 	    data_ram[  126] = 'h0000007e; 	    data_ram[  127] = 'h0000007f; 	
    data_ram[  128] = 'h00000080; 	    data_ram[  129] = 'h00000081; 	    data_ram[  130] = 'h00000082; 	    data_ram[  131] = 'h00000083; 	    data_ram[  132] = 'h00000084; 	    data_ram[  133] = 'h00000085; 	    data_ram[  134] = 'h00000086; 	    data_ram[  135] = 'h00000087; 	
    data_ram[  136] = 'h00000088; 	    data_ram[  137] = 'h00000089; 	    data_ram[  138] = 'h0000008a; 	    data_ram[  139] = 'h0000008b; 	    data_ram[  140] = 'h0000008c; 	    data_ram[  141] = 'h0000008d; 	    data_ram[  142] = 'h0000008e; 	    data_ram[  143] = 'h0000008f; 	
    data_ram[  144] = 'h00000090; 	    data_ram[  145] = 'h00000091; 	    data_ram[  146] = 'h00000092; 	    data_ram[  147] = 'h00000093; 	    data_ram[  148] = 'h00000094; 	    data_ram[  149] = 'h00000095; 	    data_ram[  150] = 'h00000096; 	    data_ram[  151] = 'h00000097; 	
    data_ram[  152] = 'h00000098; 	    data_ram[  153] = 'h00000099; 	    data_ram[  154] = 'h0000009a; 	    data_ram[  155] = 'h0000009b; 	    data_ram[  156] = 'h0000009c; 	    data_ram[  157] = 'h0000009d; 	    data_ram[  158] = 'h0000009e; 	    data_ram[  159] = 'h0000009f; 	
    data_ram[  160] = 'h000000a0; 	    data_ram[  161] = 'h000000a1; 	    data_ram[  162] = 'h000000a2; 	    data_ram[  163] = 'h000000a3; 	    data_ram[  164] = 'h000000a4; 	    data_ram[  165] = 'h000000a5; 	    data_ram[  166] = 'h000000a6; 	    data_ram[  167] = 'h000000a7; 	
    data_ram[  168] = 'h000000a8; 	    data_ram[  169] = 'h000000a9; 	    data_ram[  170] = 'h000000aa; 	    data_ram[  171] = 'h000000ab; 	    data_ram[  172] = 'h000000ac; 	    data_ram[  173] = 'h000000ad; 	    data_ram[  174] = 'h000000ae; 	    data_ram[  175] = 'h000000af; 	
    data_ram[  176] = 'h000000b0; 	    data_ram[  177] = 'h000000b1; 	    data_ram[  178] = 'h000000b2; 	    data_ram[  179] = 'h000000b3; 	    data_ram[  180] = 'h000000b4; 	    data_ram[  181] = 'h000000b5; 	    data_ram[  182] = 'h000000b6; 	    data_ram[  183] = 'h000000b7; 	
    data_ram[  184] = 'h000000b8; 	    data_ram[  185] = 'h000000b9; 	    data_ram[  186] = 'h000000ba; 	    data_ram[  187] = 'h000000bb; 	    data_ram[  188] = 'h000000bc; 	    data_ram[  189] = 'h000000bd; 	    data_ram[  190] = 'h000000be; 	    data_ram[  191] = 'h000000bf; 	
    data_ram[  192] = 'h000000c0; 	    data_ram[  193] = 'h000000c1; 	    data_ram[  194] = 'h000000c2; 	    data_ram[  195] = 'h000000c3; 	    data_ram[  196] = 'h000000c4; 	    data_ram[  197] = 'h000000c5; 	    data_ram[  198] = 'h000000c6; 	    data_ram[  199] = 'h000000c7; 	
    data_ram[  200] = 'h000000c8; 	    data_ram[  201] = 'h000000c9; 	    data_ram[  202] = 'h000000ca; 	    data_ram[  203] = 'h000000cb; 	    data_ram[  204] = 'h000000cc; 	    data_ram[  205] = 'h000000cd; 	    data_ram[  206] = 'h000000ce; 	    data_ram[  207] = 'h000000cf; 	
    data_ram[  208] = 'h000000d0; 	    data_ram[  209] = 'h000000d1; 	    data_ram[  210] = 'h000000d2; 	    data_ram[  211] = 'h000000d3; 	    data_ram[  212] = 'h000000d4; 	    data_ram[  213] = 'h000000d5; 	    data_ram[  214] = 'h000000d6; 	    data_ram[  215] = 'h000000d7; 	
    data_ram[  216] = 'h000000d8; 	    data_ram[  217] = 'h000000d9; 	    data_ram[  218] = 'h000000da; 	    data_ram[  219] = 'h000000db; 	    data_ram[  220] = 'h000000dc; 	    data_ram[  221] = 'h000000dd; 	    data_ram[  222] = 'h000000de; 	    data_ram[  223] = 'h000000df; 	
    data_ram[  224] = 'h000000e0; 	    data_ram[  225] = 'h000000e1; 	    data_ram[  226] = 'h000000e2; 	    data_ram[  227] = 'h000000e3; 	    data_ram[  228] = 'h000000e4; 	    data_ram[  229] = 'h000000e5; 	    data_ram[  230] = 'h000000e6; 	    data_ram[  231] = 'h000000e7; 	
    data_ram[  232] = 'h000000e8; 	    data_ram[  233] = 'h000000e9; 	    data_ram[  234] = 'h000000ea; 	    data_ram[  235] = 'h000000eb; 	    data_ram[  236] = 'h000000ec; 	    data_ram[  237] = 'h000000ed; 	    data_ram[  238] = 'h000000ee; 	    data_ram[  239] = 'h000000ef; 	
    data_ram[  240] = 'h000000f0; 	    data_ram[  241] = 'h000000f1; 	    data_ram[  242] = 'h000000f2; 	    data_ram[  243] = 'h000000f3; 	    data_ram[  244] = 'h000000f4; 	    data_ram[  245] = 'h000000f5; 	    data_ram[  246] = 'h000000f6; 	    data_ram[  247] = 'h000000f7; 	
    data_ram[  248] = 'h000000f8; 	    data_ram[  249] = 'h000000f9; 	    data_ram[  250] = 'h000000fa; 	    data_ram[  251] = 'h000000fb; 	    data_ram[  252] = 'h000000fc; 	    data_ram[  253] = 'h000000fd; 	    data_ram[  254] = 'h000000fe; 	    data_ram[  255] = 'h000000ff; 	
    data_ram[  256] = 'h00000100; 	    data_ram[  257] = 'h00000101; 	    data_ram[  258] = 'h00000102; 	    data_ram[  259] = 'h00000103; 	    data_ram[  260] = 'h00000104; 	    data_ram[  261] = 'h00000105; 	    data_ram[  262] = 'h00000106; 	    data_ram[  263] = 'h00000107; 	
    data_ram[  264] = 'h00000108; 	    data_ram[  265] = 'h00000109; 	    data_ram[  266] = 'h0000010a; 	    data_ram[  267] = 'h0000010b; 	    data_ram[  268] = 'h0000010c; 	    data_ram[  269] = 'h0000010d; 	    data_ram[  270] = 'h0000010e; 	    data_ram[  271] = 'h0000010f; 	
    data_ram[  272] = 'h00000110; 	    data_ram[  273] = 'h00000111; 	    data_ram[  274] = 'h00000112; 	    data_ram[  275] = 'h00000113; 	    data_ram[  276] = 'h00000114; 	    data_ram[  277] = 'h00000115; 	    data_ram[  278] = 'h00000116; 	    data_ram[  279] = 'h00000117; 	
    data_ram[  280] = 'h00000118; 	    data_ram[  281] = 'h00000119; 	    data_ram[  282] = 'h0000011a; 	    data_ram[  283] = 'h0000011b; 	    data_ram[  284] = 'h0000011c; 	    data_ram[  285] = 'h0000011d; 	    data_ram[  286] = 'h0000011e; 	    data_ram[  287] = 'h0000011f; 	
    data_ram[  288] = 'h00000120; 	    data_ram[  289] = 'h00000121; 	    data_ram[  290] = 'h00000122; 	    data_ram[  291] = 'h00000123; 	    data_ram[  292] = 'h00000124; 	    data_ram[  293] = 'h00000125; 	    data_ram[  294] = 'h00000126; 	    data_ram[  295] = 'h00000127; 	
    data_ram[  296] = 'h00000128; 	    data_ram[  297] = 'h00000129; 	    data_ram[  298] = 'h0000012a; 	    data_ram[  299] = 'h0000012b; 	    data_ram[  300] = 'h0000012c; 	    data_ram[  301] = 'h0000012d; 	    data_ram[  302] = 'h0000012e; 	    data_ram[  303] = 'h0000012f; 	
    data_ram[  304] = 'h00000130; 	    data_ram[  305] = 'h00000131; 	    data_ram[  306] = 'h00000132; 	    data_ram[  307] = 'h00000133; 	    data_ram[  308] = 'h00000134; 	    data_ram[  309] = 'h00000135; 	    data_ram[  310] = 'h00000136; 	    data_ram[  311] = 'h00000137; 	
    data_ram[  312] = 'h00000138; 	    data_ram[  313] = 'h00000139; 	    data_ram[  314] = 'h0000013a; 	    data_ram[  315] = 'h0000013b; 	    data_ram[  316] = 'h0000013c; 	    data_ram[  317] = 'h0000013d; 	    data_ram[  318] = 'h0000013e; 	    data_ram[  319] = 'h0000013f; 	
    data_ram[  320] = 'h00000140; 	    data_ram[  321] = 'h00000141; 	    data_ram[  322] = 'h00000142; 	    data_ram[  323] = 'h00000143; 	    data_ram[  324] = 'h00000144; 	    data_ram[  325] = 'h00000145; 	    data_ram[  326] = 'h00000146; 	    data_ram[  327] = 'h00000147; 	
    data_ram[  328] = 'h00000148; 	    data_ram[  329] = 'h00000149; 	    data_ram[  330] = 'h0000014a; 	    data_ram[  331] = 'h0000014b; 	    data_ram[  332] = 'h0000014c; 	    data_ram[  333] = 'h0000014d; 	    data_ram[  334] = 'h0000014e; 	    data_ram[  335] = 'h0000014f; 	
    data_ram[  336] = 'h00000150; 	    data_ram[  337] = 'h00000151; 	    data_ram[  338] = 'h00000152; 	    data_ram[  339] = 'h00000153; 	    data_ram[  340] = 'h00000154; 	    data_ram[  341] = 'h00000155; 	    data_ram[  342] = 'h00000156; 	    data_ram[  343] = 'h00000157; 	
    data_ram[  344] = 'h00000158; 	    data_ram[  345] = 'h00000159; 	    data_ram[  346] = 'h0000015a; 	    data_ram[  347] = 'h0000015b; 	    data_ram[  348] = 'h0000015c; 	    data_ram[  349] = 'h0000015d; 	    data_ram[  350] = 'h0000015e; 	    data_ram[  351] = 'h0000015f; 	
    data_ram[  352] = 'h00000160; 	    data_ram[  353] = 'h00000161; 	    data_ram[  354] = 'h00000162; 	    data_ram[  355] = 'h00000163; 	    data_ram[  356] = 'h00000164; 	    data_ram[  357] = 'h00000165; 	    data_ram[  358] = 'h00000166; 	    data_ram[  359] = 'h00000167; 	
    data_ram[  360] = 'h00000168; 	    data_ram[  361] = 'h00000169; 	    data_ram[  362] = 'h0000016a; 	    data_ram[  363] = 'h0000016b; 	    data_ram[  364] = 'h0000016c; 	    data_ram[  365] = 'h0000016d; 	    data_ram[  366] = 'h0000016e; 	    data_ram[  367] = 'h0000016f; 	
    data_ram[  368] = 'h00000170; 	    data_ram[  369] = 'h00000171; 	    data_ram[  370] = 'h00000172; 	    data_ram[  371] = 'h00000173; 	    data_ram[  372] = 'h00000174; 	    data_ram[  373] = 'h00000175; 	    data_ram[  374] = 'h00000176; 	    data_ram[  375] = 'h00000177; 	
    data_ram[  376] = 'h00000178; 	    data_ram[  377] = 'h00000179; 	    data_ram[  378] = 'h0000017a; 	    data_ram[  379] = 'h0000017b; 	    data_ram[  380] = 'h0000017c; 	    data_ram[  381] = 'h0000017d; 	    data_ram[  382] = 'h0000017e; 	    data_ram[  383] = 'h0000017f; 	
    data_ram[  384] = 'h00000180; 	    data_ram[  385] = 'h00000181; 	    data_ram[  386] = 'h00000182; 	    data_ram[  387] = 'h00000183; 	    data_ram[  388] = 'h00000184; 	    data_ram[  389] = 'h00000185; 	    data_ram[  390] = 'h00000186; 	    data_ram[  391] = 'h00000187; 	
    data_ram[  392] = 'h00000188; 	    data_ram[  393] = 'h00000189; 	    data_ram[  394] = 'h0000018a; 	    data_ram[  395] = 'h0000018b; 	    data_ram[  396] = 'h0000018c; 	    data_ram[  397] = 'h0000018d; 	    data_ram[  398] = 'h0000018e; 	    data_ram[  399] = 'h0000018f; 	
    data_ram[  400] = 'h00000190; 	    data_ram[  401] = 'h00000191; 	    data_ram[  402] = 'h00000192; 	    data_ram[  403] = 'h00000193; 	    data_ram[  404] = 'h00000194; 	    data_ram[  405] = 'h00000195; 	    data_ram[  406] = 'h00000196; 	    data_ram[  407] = 'h00000197; 	
    data_ram[  408] = 'h00000198; 	    data_ram[  409] = 'h00000199; 	    data_ram[  410] = 'h0000019a; 	    data_ram[  411] = 'h0000019b; 	    data_ram[  412] = 'h0000019c; 	    data_ram[  413] = 'h0000019d; 	    data_ram[  414] = 'h0000019e; 	    data_ram[  415] = 'h0000019f; 	
    data_ram[  416] = 'h000001a0; 	    data_ram[  417] = 'h000001a1; 	    data_ram[  418] = 'h000001a2; 	    data_ram[  419] = 'h000001a3; 	    data_ram[  420] = 'h000001a4; 	    data_ram[  421] = 'h000001a5; 	    data_ram[  422] = 'h000001a6; 	    data_ram[  423] = 'h000001a7; 	
    data_ram[  424] = 'h000001a8; 	    data_ram[  425] = 'h000001a9; 	    data_ram[  426] = 'h000001aa; 	    data_ram[  427] = 'h000001ab; 	    data_ram[  428] = 'h000001ac; 	    data_ram[  429] = 'h000001ad; 	    data_ram[  430] = 'h000001ae; 	    data_ram[  431] = 'h000001af; 	
    data_ram[  432] = 'h000001b0; 	    data_ram[  433] = 'h000001b1; 	    data_ram[  434] = 'h000001b2; 	    data_ram[  435] = 'h000001b3; 	    data_ram[  436] = 'h000001b4; 	    data_ram[  437] = 'h000001b5; 	    data_ram[  438] = 'h000001b6; 	    data_ram[  439] = 'h000001b7; 	
    data_ram[  440] = 'h000001b8; 	    data_ram[  441] = 'h000001b9; 	    data_ram[  442] = 'h000001ba; 	    data_ram[  443] = 'h000001bb; 	    data_ram[  444] = 'h000001bc; 	    data_ram[  445] = 'h000001bd; 	    data_ram[  446] = 'h000001be; 	    data_ram[  447] = 'h000001bf; 	
    data_ram[  448] = 'h000001c0; 	    data_ram[  449] = 'h000001c1; 	    data_ram[  450] = 'h000001c2; 	    data_ram[  451] = 'h000001c3; 	    data_ram[  452] = 'h000001c4; 	    data_ram[  453] = 'h000001c5; 	    data_ram[  454] = 'h000001c6; 	    data_ram[  455] = 'h000001c7; 	
    data_ram[  456] = 'h000001c8; 	    data_ram[  457] = 'h000001c9; 	    data_ram[  458] = 'h000001ca; 	    data_ram[  459] = 'h000001cb; 	    data_ram[  460] = 'h000001cc; 	    data_ram[  461] = 'h000001cd; 	    data_ram[  462] = 'h000001ce; 	    data_ram[  463] = 'h000001cf; 	
    data_ram[  464] = 'h000001d0; 	    data_ram[  465] = 'h000001d1; 	    data_ram[  466] = 'h000001d2; 	    data_ram[  467] = 'h000001d3; 	    data_ram[  468] = 'h000001d4; 	    data_ram[  469] = 'h000001d5; 	    data_ram[  470] = 'h000001d6; 	    data_ram[  471] = 'h000001d7; 	
    data_ram[  472] = 'h000001d8; 	    data_ram[  473] = 'h000001d9; 	    data_ram[  474] = 'h000001da; 	    data_ram[  475] = 'h000001db; 	    data_ram[  476] = 'h000001dc; 	    data_ram[  477] = 'h000001dd; 	    data_ram[  478] = 'h000001de; 	    data_ram[  479] = 'h000001df; 	
    data_ram[  480] = 'h000001e0; 	    data_ram[  481] = 'h000001e1; 	    data_ram[  482] = 'h000001e2; 	    data_ram[  483] = 'h000001e3; 	    data_ram[  484] = 'h000001e4; 	    data_ram[  485] = 'h000001e5; 	    data_ram[  486] = 'h000001e6; 	    data_ram[  487] = 'h000001e7; 	
    data_ram[  488] = 'h000001e8; 	    data_ram[  489] = 'h000001e9; 	    data_ram[  490] = 'h000001ea; 	    data_ram[  491] = 'h000001eb; 	    data_ram[  492] = 'h000001ec; 	    data_ram[  493] = 'h000001ed; 	    data_ram[  494] = 'h000001ee; 	    data_ram[  495] = 'h000001ef; 	
    data_ram[  496] = 'h000001f0; 	    data_ram[  497] = 'h000001f1; 	    data_ram[  498] = 'h000001f2; 	    data_ram[  499] = 'h000001f3; 	    data_ram[  500] = 'h000001f4; 	    data_ram[  501] = 'h000001f5; 	    data_ram[  502] = 'h000001f6; 	    data_ram[  503] = 'h000001f7; 	
    data_ram[  504] = 'h000001f8; 	    data_ram[  505] = 'h000001f9; 	    data_ram[  506] = 'h000001fa; 	    data_ram[  507] = 'h000001fb; 	    data_ram[  508] = 'h000001fc; 	    data_ram[  509] = 'h000001fd; 	    data_ram[  510] = 'h000001fe; 	    data_ram[  511] = 'h000001ff; 	
    data_ram[  512] = 'h00000200; 	    data_ram[  513] = 'h00000201; 	    data_ram[  514] = 'h00000202; 	    data_ram[  515] = 'h00000203; 	    data_ram[  516] = 'h00000204; 	    data_ram[  517] = 'h00000205; 	    data_ram[  518] = 'h00000206; 	    data_ram[  519] = 'h00000207; 	
    data_ram[  520] = 'h00000208; 	    data_ram[  521] = 'h00000209; 	    data_ram[  522] = 'h0000020a; 	    data_ram[  523] = 'h0000020b; 	    data_ram[  524] = 'h0000020c; 	    data_ram[  525] = 'h0000020d; 	    data_ram[  526] = 'h0000020e; 	    data_ram[  527] = 'h0000020f; 	
    data_ram[  528] = 'h00000210; 	    data_ram[  529] = 'h00000211; 	    data_ram[  530] = 'h00000212; 	    data_ram[  531] = 'h00000213; 	    data_ram[  532] = 'h00000214; 	    data_ram[  533] = 'h00000215; 	    data_ram[  534] = 'h00000216; 	    data_ram[  535] = 'h00000217; 	
    data_ram[  536] = 'h00000218; 	    data_ram[  537] = 'h00000219; 	    data_ram[  538] = 'h0000021a; 	    data_ram[  539] = 'h0000021b; 	    data_ram[  540] = 'h0000021c; 	    data_ram[  541] = 'h0000021d; 	    data_ram[  542] = 'h0000021e; 	    data_ram[  543] = 'h0000021f; 	
    data_ram[  544] = 'h00000220; 	    data_ram[  545] = 'h00000221; 	    data_ram[  546] = 'h00000222; 	    data_ram[  547] = 'h00000223; 	    data_ram[  548] = 'h00000224; 	    data_ram[  549] = 'h00000225; 	    data_ram[  550] = 'h00000226; 	    data_ram[  551] = 'h00000227; 	
    data_ram[  552] = 'h00000228; 	    data_ram[  553] = 'h00000229; 	    data_ram[  554] = 'h0000022a; 	    data_ram[  555] = 'h0000022b; 	    data_ram[  556] = 'h0000022c; 	    data_ram[  557] = 'h0000022d; 	    data_ram[  558] = 'h0000022e; 	    data_ram[  559] = 'h0000022f; 	
    data_ram[  560] = 'h00000230; 	    data_ram[  561] = 'h00000231; 	    data_ram[  562] = 'h00000232; 	    data_ram[  563] = 'h00000233; 	    data_ram[  564] = 'h00000234; 	    data_ram[  565] = 'h00000235; 	    data_ram[  566] = 'h00000236; 	    data_ram[  567] = 'h00000237; 	
    data_ram[  568] = 'h00000238; 	    data_ram[  569] = 'h00000239; 	    data_ram[  570] = 'h0000023a; 	    data_ram[  571] = 'h0000023b; 	    data_ram[  572] = 'h0000023c; 	    data_ram[  573] = 'h0000023d; 	    data_ram[  574] = 'h0000023e; 	    data_ram[  575] = 'h0000023f; 	
    data_ram[  576] = 'h00000240; 	    data_ram[  577] = 'h00000241; 	    data_ram[  578] = 'h00000242; 	    data_ram[  579] = 'h00000243; 	    data_ram[  580] = 'h00000244; 	    data_ram[  581] = 'h00000245; 	    data_ram[  582] = 'h00000246; 	    data_ram[  583] = 'h00000247; 	
    data_ram[  584] = 'h00000248; 	    data_ram[  585] = 'h00000249; 	    data_ram[  586] = 'h0000024a; 	    data_ram[  587] = 'h0000024b; 	    data_ram[  588] = 'h0000024c; 	    data_ram[  589] = 'h0000024d; 	    data_ram[  590] = 'h0000024e; 	    data_ram[  591] = 'h0000024f; 	
    data_ram[  592] = 'h00000250; 	    data_ram[  593] = 'h00000251; 	    data_ram[  594] = 'h00000252; 	    data_ram[  595] = 'h00000253; 	    data_ram[  596] = 'h00000254; 	    data_ram[  597] = 'h00000255; 	    data_ram[  598] = 'h00000256; 	    data_ram[  599] = 'h00000257; 	
    data_ram[  600] = 'h00000258; 	    data_ram[  601] = 'h00000259; 	    data_ram[  602] = 'h0000025a; 	    data_ram[  603] = 'h0000025b; 	    data_ram[  604] = 'h0000025c; 	    data_ram[  605] = 'h0000025d; 	    data_ram[  606] = 'h0000025e; 	    data_ram[  607] = 'h0000025f; 	
    data_ram[  608] = 'h00000260; 	    data_ram[  609] = 'h00000261; 	    data_ram[  610] = 'h00000262; 	    data_ram[  611] = 'h00000263; 	    data_ram[  612] = 'h00000264; 	    data_ram[  613] = 'h00000265; 	    data_ram[  614] = 'h00000266; 	    data_ram[  615] = 'h00000267; 	
    data_ram[  616] = 'h00000268; 	    data_ram[  617] = 'h00000269; 	    data_ram[  618] = 'h0000026a; 	    data_ram[  619] = 'h0000026b; 	    data_ram[  620] = 'h0000026c; 	    data_ram[  621] = 'h0000026d; 	    data_ram[  622] = 'h0000026e; 	    data_ram[  623] = 'h0000026f; 	
    data_ram[  624] = 'h00000270; 	    data_ram[  625] = 'h00000271; 	    data_ram[  626] = 'h00000272; 	    data_ram[  627] = 'h00000273; 	    data_ram[  628] = 'h00000274; 	    data_ram[  629] = 'h00000275; 	    data_ram[  630] = 'h00000276; 	    data_ram[  631] = 'h00000277; 	
    data_ram[  632] = 'h00000278; 	    data_ram[  633] = 'h00000279; 	    data_ram[  634] = 'h0000027a; 	    data_ram[  635] = 'h0000027b; 	    data_ram[  636] = 'h0000027c; 	    data_ram[  637] = 'h0000027d; 	    data_ram[  638] = 'h0000027e; 	    data_ram[  639] = 'h0000027f; 	
    data_ram[  640] = 'h00000280; 	    data_ram[  641] = 'h00000281; 	    data_ram[  642] = 'h00000282; 	    data_ram[  643] = 'h00000283; 	    data_ram[  644] = 'h00000284; 	    data_ram[  645] = 'h00000285; 	    data_ram[  646] = 'h00000286; 	    data_ram[  647] = 'h00000287; 	
    data_ram[  648] = 'h00000288; 	    data_ram[  649] = 'h00000289; 	    data_ram[  650] = 'h0000028a; 	    data_ram[  651] = 'h0000028b; 	    data_ram[  652] = 'h0000028c; 	    data_ram[  653] = 'h0000028d; 	    data_ram[  654] = 'h0000028e; 	    data_ram[  655] = 'h0000028f; 	
    data_ram[  656] = 'h00000290; 	    data_ram[  657] = 'h00000291; 	    data_ram[  658] = 'h00000292; 	    data_ram[  659] = 'h00000293; 	    data_ram[  660] = 'h00000294; 	    data_ram[  661] = 'h00000295; 	    data_ram[  662] = 'h00000296; 	    data_ram[  663] = 'h00000297; 	
    data_ram[  664] = 'h00000298; 	    data_ram[  665] = 'h00000299; 	    data_ram[  666] = 'h0000029a; 	    data_ram[  667] = 'h0000029b; 	    data_ram[  668] = 'h0000029c; 	    data_ram[  669] = 'h0000029d; 	    data_ram[  670] = 'h0000029e; 	    data_ram[  671] = 'h0000029f; 	
    data_ram[  672] = 'h000002a0; 	    data_ram[  673] = 'h000002a1; 	    data_ram[  674] = 'h000002a2; 	    data_ram[  675] = 'h000002a3; 	    data_ram[  676] = 'h000002a4; 	    data_ram[  677] = 'h000002a5; 	    data_ram[  678] = 'h000002a6; 	    data_ram[  679] = 'h000002a7; 	
    data_ram[  680] = 'h000002a8; 	    data_ram[  681] = 'h000002a9; 	    data_ram[  682] = 'h000002aa; 	    data_ram[  683] = 'h000002ab; 	    data_ram[  684] = 'h000002ac; 	    data_ram[  685] = 'h000002ad; 	    data_ram[  686] = 'h000002ae; 	    data_ram[  687] = 'h000002af; 	
    data_ram[  688] = 'h000002b0; 	    data_ram[  689] = 'h000002b1; 	    data_ram[  690] = 'h000002b2; 	    data_ram[  691] = 'h000002b3; 	    data_ram[  692] = 'h000002b4; 	    data_ram[  693] = 'h000002b5; 	    data_ram[  694] = 'h000002b6; 	    data_ram[  695] = 'h000002b7; 	
    data_ram[  696] = 'h000002b8; 	    data_ram[  697] = 'h000002b9; 	    data_ram[  698] = 'h000002ba; 	    data_ram[  699] = 'h000002bb; 	    data_ram[  700] = 'h000002bc; 	    data_ram[  701] = 'h000002bd; 	    data_ram[  702] = 'h000002be; 	    data_ram[  703] = 'h000002bf; 	
    data_ram[  704] = 'h000002c0; 	    data_ram[  705] = 'h000002c1; 	    data_ram[  706] = 'h000002c2; 	    data_ram[  707] = 'h000002c3; 	    data_ram[  708] = 'h000002c4; 	    data_ram[  709] = 'h000002c5; 	    data_ram[  710] = 'h000002c6; 	    data_ram[  711] = 'h000002c7; 	
    data_ram[  712] = 'h000002c8; 	    data_ram[  713] = 'h000002c9; 	    data_ram[  714] = 'h000002ca; 	    data_ram[  715] = 'h000002cb; 	    data_ram[  716] = 'h000002cc; 	    data_ram[  717] = 'h000002cd; 	    data_ram[  718] = 'h000002ce; 	    data_ram[  719] = 'h000002cf; 	
    data_ram[  720] = 'h000002d0; 	    data_ram[  721] = 'h000002d1; 	    data_ram[  722] = 'h000002d2; 	    data_ram[  723] = 'h000002d3; 	    data_ram[  724] = 'h000002d4; 	    data_ram[  725] = 'h000002d5; 	    data_ram[  726] = 'h000002d6; 	    data_ram[  727] = 'h000002d7; 	
    data_ram[  728] = 'h000002d8; 	    data_ram[  729] = 'h000002d9; 	    data_ram[  730] = 'h000002da; 	    data_ram[  731] = 'h000002db; 	    data_ram[  732] = 'h000002dc; 	    data_ram[  733] = 'h000002dd; 	    data_ram[  734] = 'h000002de; 	    data_ram[  735] = 'h000002df; 	
    data_ram[  736] = 'h000002e0; 	    data_ram[  737] = 'h000002e1; 	    data_ram[  738] = 'h000002e2; 	    data_ram[  739] = 'h000002e3; 	    data_ram[  740] = 'h000002e4; 	    data_ram[  741] = 'h000002e5; 	    data_ram[  742] = 'h000002e6; 	    data_ram[  743] = 'h000002e7; 	
    data_ram[  744] = 'h000002e8; 	    data_ram[  745] = 'h000002e9; 	    data_ram[  746] = 'h000002ea; 	    data_ram[  747] = 'h000002eb; 	    data_ram[  748] = 'h000002ec; 	    data_ram[  749] = 'h000002ed; 	    data_ram[  750] = 'h000002ee; 	    data_ram[  751] = 'h000002ef; 	
    data_ram[  752] = 'h000002f0; 	    data_ram[  753] = 'h000002f1; 	    data_ram[  754] = 'h000002f2; 	    data_ram[  755] = 'h000002f3; 	    data_ram[  756] = 'h000002f4; 	    data_ram[  757] = 'h000002f5; 	    data_ram[  758] = 'h000002f6; 	    data_ram[  759] = 'h000002f7; 	
    data_ram[  760] = 'h000002f8; 	    data_ram[  761] = 'h000002f9; 	    data_ram[  762] = 'h000002fa; 	    data_ram[  763] = 'h000002fb; 	    data_ram[  764] = 'h000002fc; 	    data_ram[  765] = 'h000002fd; 	    data_ram[  766] = 'h000002fe; 	    data_ram[  767] = 'h000002ff; 	
    data_ram[  768] = 'h00000300; 	    data_ram[  769] = 'h00000301; 	    data_ram[  770] = 'h00000302; 	    data_ram[  771] = 'h00000303; 	    data_ram[  772] = 'h00000304; 	    data_ram[  773] = 'h00000305; 	    data_ram[  774] = 'h00000306; 	    data_ram[  775] = 'h00000307; 	
    data_ram[  776] = 'h00000308; 	    data_ram[  777] = 'h00000309; 	    data_ram[  778] = 'h0000030a; 	    data_ram[  779] = 'h0000030b; 	    data_ram[  780] = 'h0000030c; 	    data_ram[  781] = 'h0000030d; 	    data_ram[  782] = 'h0000030e; 	    data_ram[  783] = 'h0000030f; 	
    data_ram[  784] = 'h00000310; 	    data_ram[  785] = 'h00000311; 	    data_ram[  786] = 'h00000312; 	    data_ram[  787] = 'h00000313; 	    data_ram[  788] = 'h00000314; 	    data_ram[  789] = 'h00000315; 	    data_ram[  790] = 'h00000316; 	    data_ram[  791] = 'h00000317; 	
    data_ram[  792] = 'h00000318; 	    data_ram[  793] = 'h00000319; 	    data_ram[  794] = 'h0000031a; 	    data_ram[  795] = 'h0000031b; 	    data_ram[  796] = 'h0000031c; 	    data_ram[  797] = 'h0000031d; 	    data_ram[  798] = 'h0000031e; 	    data_ram[  799] = 'h0000031f; 	
    data_ram[  800] = 'h00000320; 	    data_ram[  801] = 'h00000321; 	    data_ram[  802] = 'h00000322; 	    data_ram[  803] = 'h00000323; 	    data_ram[  804] = 'h00000324; 	    data_ram[  805] = 'h00000325; 	    data_ram[  806] = 'h00000326; 	    data_ram[  807] = 'h00000327; 	
    data_ram[  808] = 'h00000328; 	    data_ram[  809] = 'h00000329; 	    data_ram[  810] = 'h0000032a; 	    data_ram[  811] = 'h0000032b; 	    data_ram[  812] = 'h0000032c; 	    data_ram[  813] = 'h0000032d; 	    data_ram[  814] = 'h0000032e; 	    data_ram[  815] = 'h0000032f; 	
    data_ram[  816] = 'h00000330; 	    data_ram[  817] = 'h00000331; 	    data_ram[  818] = 'h00000332; 	    data_ram[  819] = 'h00000333; 	    data_ram[  820] = 'h00000334; 	    data_ram[  821] = 'h00000335; 	    data_ram[  822] = 'h00000336; 	    data_ram[  823] = 'h00000337; 	
    data_ram[  824] = 'h00000338; 	    data_ram[  825] = 'h00000339; 	    data_ram[  826] = 'h0000033a; 	    data_ram[  827] = 'h0000033b; 	    data_ram[  828] = 'h0000033c; 	    data_ram[  829] = 'h0000033d; 	    data_ram[  830] = 'h0000033e; 	    data_ram[  831] = 'h0000033f; 	
    data_ram[  832] = 'h00000340; 	    data_ram[  833] = 'h00000341; 	    data_ram[  834] = 'h00000342; 	    data_ram[  835] = 'h00000343; 	    data_ram[  836] = 'h00000344; 	    data_ram[  837] = 'h00000345; 	    data_ram[  838] = 'h00000346; 	    data_ram[  839] = 'h00000347; 	
    data_ram[  840] = 'h00000348; 	    data_ram[  841] = 'h00000349; 	    data_ram[  842] = 'h0000034a; 	    data_ram[  843] = 'h0000034b; 	    data_ram[  844] = 'h0000034c; 	    data_ram[  845] = 'h0000034d; 	    data_ram[  846] = 'h0000034e; 	    data_ram[  847] = 'h0000034f; 	
    data_ram[  848] = 'h00000350; 	    data_ram[  849] = 'h00000351; 	    data_ram[  850] = 'h00000352; 	    data_ram[  851] = 'h00000353; 	    data_ram[  852] = 'h00000354; 	    data_ram[  853] = 'h00000355; 	    data_ram[  854] = 'h00000356; 	    data_ram[  855] = 'h00000357; 	
    data_ram[  856] = 'h00000358; 	    data_ram[  857] = 'h00000359; 	    data_ram[  858] = 'h0000035a; 	    data_ram[  859] = 'h0000035b; 	    data_ram[  860] = 'h0000035c; 	    data_ram[  861] = 'h0000035d; 	    data_ram[  862] = 'h0000035e; 	    data_ram[  863] = 'h0000035f; 	
    data_ram[  864] = 'h00000360; 	    data_ram[  865] = 'h00000361; 	    data_ram[  866] = 'h00000362; 	    data_ram[  867] = 'h00000363; 	    data_ram[  868] = 'h00000364; 	    data_ram[  869] = 'h00000365; 	    data_ram[  870] = 'h00000366; 	    data_ram[  871] = 'h00000367; 	
    data_ram[  872] = 'h00000368; 	    data_ram[  873] = 'h00000369; 	    data_ram[  874] = 'h0000036a; 	    data_ram[  875] = 'h0000036b; 	    data_ram[  876] = 'h0000036c; 	    data_ram[  877] = 'h0000036d; 	    data_ram[  878] = 'h0000036e; 	    data_ram[  879] = 'h0000036f; 	
    data_ram[  880] = 'h00000370; 	    data_ram[  881] = 'h00000371; 	    data_ram[  882] = 'h00000372; 	    data_ram[  883] = 'h00000373; 	    data_ram[  884] = 'h00000374; 	    data_ram[  885] = 'h00000375; 	    data_ram[  886] = 'h00000376; 	    data_ram[  887] = 'h00000377; 	
    data_ram[  888] = 'h00000378; 	    data_ram[  889] = 'h00000379; 	    data_ram[  890] = 'h0000037a; 	    data_ram[  891] = 'h0000037b; 	    data_ram[  892] = 'h0000037c; 	    data_ram[  893] = 'h0000037d; 	    data_ram[  894] = 'h0000037e; 	    data_ram[  895] = 'h0000037f; 	
    data_ram[  896] = 'h00000380; 	    data_ram[  897] = 'h00000381; 	    data_ram[  898] = 'h00000382; 	    data_ram[  899] = 'h00000383; 	    data_ram[  900] = 'h00000384; 	    data_ram[  901] = 'h00000385; 	    data_ram[  902] = 'h00000386; 	    data_ram[  903] = 'h00000387; 	
    data_ram[  904] = 'h00000388; 	    data_ram[  905] = 'h00000389; 	    data_ram[  906] = 'h0000038a; 	    data_ram[  907] = 'h0000038b; 	    data_ram[  908] = 'h0000038c; 	    data_ram[  909] = 'h0000038d; 	    data_ram[  910] = 'h0000038e; 	    data_ram[  911] = 'h0000038f; 	
    data_ram[  912] = 'h00000390; 	    data_ram[  913] = 'h00000391; 	    data_ram[  914] = 'h00000392; 	    data_ram[  915] = 'h00000393; 	    data_ram[  916] = 'h00000394; 	    data_ram[  917] = 'h00000395; 	    data_ram[  918] = 'h00000396; 	    data_ram[  919] = 'h00000397; 	
    data_ram[  920] = 'h00000398; 	    data_ram[  921] = 'h00000399; 	    data_ram[  922] = 'h0000039a; 	    data_ram[  923] = 'h0000039b; 	    data_ram[  924] = 'h0000039c; 	    data_ram[  925] = 'h0000039d; 	    data_ram[  926] = 'h0000039e; 	    data_ram[  927] = 'h0000039f; 	
    data_ram[  928] = 'h000003a0; 	    data_ram[  929] = 'h000003a1; 	    data_ram[  930] = 'h000003a2; 	    data_ram[  931] = 'h000003a3; 	    data_ram[  932] = 'h000003a4; 	    data_ram[  933] = 'h000003a5; 	    data_ram[  934] = 'h000003a6; 	    data_ram[  935] = 'h000003a7; 	
    data_ram[  936] = 'h000003a8; 	    data_ram[  937] = 'h000003a9; 	    data_ram[  938] = 'h000003aa; 	    data_ram[  939] = 'h000003ab; 	    data_ram[  940] = 'h000003ac; 	    data_ram[  941] = 'h000003ad; 	    data_ram[  942] = 'h000003ae; 	    data_ram[  943] = 'h000003af; 	
    data_ram[  944] = 'h000003b0; 	    data_ram[  945] = 'h000003b1; 	    data_ram[  946] = 'h000003b2; 	    data_ram[  947] = 'h000003b3; 	    data_ram[  948] = 'h000003b4; 	    data_ram[  949] = 'h000003b5; 	    data_ram[  950] = 'h000003b6; 	    data_ram[  951] = 'h000003b7; 	
    data_ram[  952] = 'h000003b8; 	    data_ram[  953] = 'h000003b9; 	    data_ram[  954] = 'h000003ba; 	    data_ram[  955] = 'h000003bb; 	    data_ram[  956] = 'h000003bc; 	    data_ram[  957] = 'h000003bd; 	    data_ram[  958] = 'h000003be; 	    data_ram[  959] = 'h000003bf; 	
    data_ram[  960] = 'h000003c0; 	    data_ram[  961] = 'h000003c1; 	    data_ram[  962] = 'h000003c2; 	    data_ram[  963] = 'h000003c3; 	    data_ram[  964] = 'h000003c4; 	    data_ram[  965] = 'h000003c5; 	    data_ram[  966] = 'h000003c6; 	    data_ram[  967] = 'h000003c7; 	
    data_ram[  968] = 'h000003c8; 	    data_ram[  969] = 'h000003c9; 	    data_ram[  970] = 'h000003ca; 	    data_ram[  971] = 'h000003cb; 	    data_ram[  972] = 'h000003cc; 	    data_ram[  973] = 'h000003cd; 	    data_ram[  974] = 'h000003ce; 	    data_ram[  975] = 'h000003cf; 	
    data_ram[  976] = 'h000003d0; 	    data_ram[  977] = 'h000003d1; 	    data_ram[  978] = 'h000003d2; 	    data_ram[  979] = 'h000003d3; 	    data_ram[  980] = 'h000003d4; 	    data_ram[  981] = 'h000003d5; 	    data_ram[  982] = 'h000003d6; 	    data_ram[  983] = 'h000003d7; 	
    data_ram[  984] = 'h000003d8; 	    data_ram[  985] = 'h000003d9; 	    data_ram[  986] = 'h000003da; 	    data_ram[  987] = 'h000003db; 	    data_ram[  988] = 'h000003dc; 	    data_ram[  989] = 'h000003dd; 	    data_ram[  990] = 'h000003de; 	    data_ram[  991] = 'h000003df; 	
    data_ram[  992] = 'h000003e0; 	    data_ram[  993] = 'h000003e1; 	    data_ram[  994] = 'h000003e2; 	    data_ram[  995] = 'h000003e3; 	    data_ram[  996] = 'h000003e4; 	    data_ram[  997] = 'h000003e5; 	    data_ram[  998] = 'h000003e6; 	    data_ram[  999] = 'h000003e7; 	
    data_ram[ 1000] = 'h000003e8; 	    data_ram[ 1001] = 'h000003e9; 	    data_ram[ 1002] = 'h000003ea; 	    data_ram[ 1003] = 'h000003eb; 	    data_ram[ 1004] = 'h000003ec; 	    data_ram[ 1005] = 'h000003ed; 	    data_ram[ 1006] = 'h000003ee; 	    data_ram[ 1007] = 'h000003ef; 	
    data_ram[ 1008] = 'h000003f0; 	    data_ram[ 1009] = 'h000003f1; 	    data_ram[ 1010] = 'h000003f2; 	    data_ram[ 1011] = 'h000003f3; 	    data_ram[ 1012] = 'h000003f4; 	    data_ram[ 1013] = 'h000003f5; 	    data_ram[ 1014] = 'h000003f6; 	    data_ram[ 1015] = 'h000003f7; 	
    data_ram[ 1016] = 'h000003f8; 	    data_ram[ 1017] = 'h000003f9; 	    data_ram[ 1018] = 'h000003fa; 	    data_ram[ 1019] = 'h000003fb; 	    data_ram[ 1020] = 'h000003fc; 	    data_ram[ 1021] = 'h000003fd; 	    data_ram[ 1022] = 'h000003fe; 	    data_ram[ 1023] = 'h000003ff; 	

end
initial begin
    i_addr_rom[    0] = 'h000001b0; 	    d_addr_rom[    0] = 'h00000eac; 	    wdata_rom[    0] = 'hbbbbea4a; 	    wvalid_rom[    0] = 0; 
    i_addr_rom[    1] = 'h000000ac; 	    d_addr_rom[    1] = 'h00000810; 	    wdata_rom[    1] = 'h89c9f387; 	    wvalid_rom[    1] = 0; 
    i_addr_rom[    2] = 'h00000538; 	    d_addr_rom[    2] = 'h0000098c; 	    wdata_rom[    2] = 'h89375bd2; 	    wvalid_rom[    2] = 1; 
    i_addr_rom[    3] = 'h00000478; 	    d_addr_rom[    3] = 'h000009e8; 	    wdata_rom[    3] = 'h865cbbd8; 	    wvalid_rom[    3] = 1; 
    i_addr_rom[    4] = 'h000002c4; 	    d_addr_rom[    4] = 'h00000ac8; 	    wdata_rom[    4] = 'h644bf05e; 	    wvalid_rom[    4] = 0; 
    i_addr_rom[    5] = 'h00000664; 	    d_addr_rom[    5] = 'h00000c6c; 	    wdata_rom[    5] = 'hccaf697d; 	    wvalid_rom[    5] = 0; 
    i_addr_rom[    6] = 'h00000598; 	    d_addr_rom[    6] = 'h00000c0c; 	    wdata_rom[    6] = 'h660d4262; 	    wvalid_rom[    6] = 1; 
    i_addr_rom[    7] = 'h0000066c; 	    d_addr_rom[    7] = 'h00000bb4; 	    wdata_rom[    7] = 'hd8b9db33; 	    wvalid_rom[    7] = 0; 
    i_addr_rom[    8] = 'h00000220; 	    d_addr_rom[    8] = 'h00000814; 	    wdata_rom[    8] = 'hc95993ea; 	    wvalid_rom[    8] = 0; 
    i_addr_rom[    9] = 'h000007d8; 	    d_addr_rom[    9] = 'h00000cf8; 	    wdata_rom[    9] = 'h7e8ef0d1; 	    wvalid_rom[    9] = 1; 
    i_addr_rom[   10] = 'h00000454; 	    d_addr_rom[   10] = 'h00000f28; 	    wdata_rom[   10] = 'hc9c9e412; 	    wvalid_rom[   10] = 1; 
    i_addr_rom[   11] = 'h00000270; 	    d_addr_rom[   11] = 'h00000c4c; 	    wdata_rom[   11] = 'hcf33d4ba; 	    wvalid_rom[   11] = 1; 
    i_addr_rom[   12] = 'h00000134; 	    d_addr_rom[   12] = 'h00000888; 	    wdata_rom[   12] = 'h53aa623e; 	    wvalid_rom[   12] = 1; 
    i_addr_rom[   13] = 'h00000114; 	    d_addr_rom[   13] = 'h00000844; 	    wdata_rom[   13] = 'hd4e694e1; 	    wvalid_rom[   13] = 1; 
    i_addr_rom[   14] = 'h00000604; 	    d_addr_rom[   14] = 'h00000fe0; 	    wdata_rom[   14] = 'hb2aee417; 	    wvalid_rom[   14] = 1; 
    i_addr_rom[   15] = 'h000004ec; 	    d_addr_rom[   15] = 'h0000094c; 	    wdata_rom[   15] = 'h22b71ca3; 	    wvalid_rom[   15] = 0; 
    i_addr_rom[   16] = 'h0000031c; 	    d_addr_rom[   16] = 'h000008b4; 	    wdata_rom[   16] = 'hd8653a11; 	    wvalid_rom[   16] = 0; 
    i_addr_rom[   17] = 'h0000012c; 	    d_addr_rom[   17] = 'h00000820; 	    wdata_rom[   17] = 'he074a661; 	    wvalid_rom[   17] = 1; 
    i_addr_rom[   18] = 'h00000098; 	    d_addr_rom[   18] = 'h00000800; 	    wdata_rom[   18] = 'h1513bf12; 	    wvalid_rom[   18] = 0; 
    i_addr_rom[   19] = 'h000004c0; 	    d_addr_rom[   19] = 'h00000c8c; 	    wdata_rom[   19] = 'he02500a3; 	    wvalid_rom[   19] = 0; 
    i_addr_rom[   20] = 'h000001d4; 	    d_addr_rom[   20] = 'h00000cec; 	    wdata_rom[   20] = 'hc8f0e9c1; 	    wvalid_rom[   20] = 1; 
    i_addr_rom[   21] = 'h00000494; 	    d_addr_rom[   21] = 'h00000a80; 	    wdata_rom[   21] = 'h1bc24f00; 	    wvalid_rom[   21] = 1; 
    i_addr_rom[   22] = 'h00000738; 	    d_addr_rom[   22] = 'h00000940; 	    wdata_rom[   22] = 'h777e05a2; 	    wvalid_rom[   22] = 1; 
    i_addr_rom[   23] = 'h00000138; 	    d_addr_rom[   23] = 'h00000f58; 	    wdata_rom[   23] = 'h0348268e; 	    wvalid_rom[   23] = 1; 
    i_addr_rom[   24] = 'h00000208; 	    d_addr_rom[   24] = 'h00000cfc; 	    wdata_rom[   24] = 'haee03ecd; 	    wvalid_rom[   24] = 1; 
    i_addr_rom[   25] = 'h000000d8; 	    d_addr_rom[   25] = 'h00000c7c; 	    wdata_rom[   25] = 'hdb038347; 	    wvalid_rom[   25] = 0; 
    i_addr_rom[   26] = 'h000004fc; 	    d_addr_rom[   26] = 'h00000e6c; 	    wdata_rom[   26] = 'he42b413b; 	    wvalid_rom[   26] = 1; 
    i_addr_rom[   27] = 'h0000011c; 	    d_addr_rom[   27] = 'h00000e64; 	    wdata_rom[   27] = 'h33dd9c8b; 	    wvalid_rom[   27] = 1; 
    i_addr_rom[   28] = 'h00000780; 	    d_addr_rom[   28] = 'h00000eb4; 	    wdata_rom[   28] = 'hc53c8a3e; 	    wvalid_rom[   28] = 0; 
    i_addr_rom[   29] = 'h000004b4; 	    d_addr_rom[   29] = 'h00000eac; 	    wdata_rom[   29] = 'h54e10299; 	    wvalid_rom[   29] = 0; 
    i_addr_rom[   30] = 'h00000340; 	    d_addr_rom[   30] = 'h00000f0c; 	    wdata_rom[   30] = 'h3922c286; 	    wvalid_rom[   30] = 1; 
    i_addr_rom[   31] = 'h00000198; 	    d_addr_rom[   31] = 'h00000834; 	    wdata_rom[   31] = 'h0e108b7c; 	    wvalid_rom[   31] = 0; 
    i_addr_rom[   32] = 'h00000264; 	    d_addr_rom[   32] = 'h0000095c; 	    wdata_rom[   32] = 'hc778abe4; 	    wvalid_rom[   32] = 1; 
    i_addr_rom[   33] = 'h00000410; 	    d_addr_rom[   33] = 'h00000988; 	    wdata_rom[   33] = 'hed2140ac; 	    wvalid_rom[   33] = 1; 
    i_addr_rom[   34] = 'h00000358; 	    d_addr_rom[   34] = 'h0000086c; 	    wdata_rom[   34] = 'h55babd53; 	    wvalid_rom[   34] = 1; 
    i_addr_rom[   35] = 'h000006f8; 	    d_addr_rom[   35] = 'h00000abc; 	    wdata_rom[   35] = 'h63af23c8; 	    wvalid_rom[   35] = 1; 
    i_addr_rom[   36] = 'h0000050c; 	    d_addr_rom[   36] = 'h000008a4; 	    wdata_rom[   36] = 'hcaa02e5c; 	    wvalid_rom[   36] = 1; 
    i_addr_rom[   37] = 'h00000234; 	    d_addr_rom[   37] = 'h00000b00; 	    wdata_rom[   37] = 'hffcda3ff; 	    wvalid_rom[   37] = 0; 
    i_addr_rom[   38] = 'h000006c0; 	    d_addr_rom[   38] = 'h00000850; 	    wdata_rom[   38] = 'he561fdd9; 	    wvalid_rom[   38] = 0; 
    i_addr_rom[   39] = 'h00000170; 	    d_addr_rom[   39] = 'h00000f70; 	    wdata_rom[   39] = 'h70f28b65; 	    wvalid_rom[   39] = 0; 
    i_addr_rom[   40] = 'h000000a4; 	    d_addr_rom[   40] = 'h00000cf0; 	    wdata_rom[   40] = 'hc50849b3; 	    wvalid_rom[   40] = 1; 
    i_addr_rom[   41] = 'h00000284; 	    d_addr_rom[   41] = 'h00000d0c; 	    wdata_rom[   41] = 'h4e44658a; 	    wvalid_rom[   41] = 0; 
    i_addr_rom[   42] = 'h000002ac; 	    d_addr_rom[   42] = 'h000009cc; 	    wdata_rom[   42] = 'hc627712e; 	    wvalid_rom[   42] = 0; 
    i_addr_rom[   43] = 'h00000290; 	    d_addr_rom[   43] = 'h00000f30; 	    wdata_rom[   43] = 'h33a0092a; 	    wvalid_rom[   43] = 1; 
    i_addr_rom[   44] = 'h000003a8; 	    d_addr_rom[   44] = 'h00000e2c; 	    wdata_rom[   44] = 'he75d8844; 	    wvalid_rom[   44] = 1; 
    i_addr_rom[   45] = 'h000007dc; 	    d_addr_rom[   45] = 'h00000ab4; 	    wdata_rom[   45] = 'h3bb91b55; 	    wvalid_rom[   45] = 1; 
    i_addr_rom[   46] = 'h0000024c; 	    d_addr_rom[   46] = 'h00000ab0; 	    wdata_rom[   46] = 'hfd66956a; 	    wvalid_rom[   46] = 1; 
    i_addr_rom[   47] = 'h000000b4; 	    d_addr_rom[   47] = 'h00000848; 	    wdata_rom[   47] = 'h9ea88fb2; 	    wvalid_rom[   47] = 0; 
    i_addr_rom[   48] = 'h000001f4; 	    d_addr_rom[   48] = 'h0000087c; 	    wdata_rom[   48] = 'h04c771bf; 	    wvalid_rom[   48] = 1; 
    i_addr_rom[   49] = 'h00000278; 	    d_addr_rom[   49] = 'h0000098c; 	    wdata_rom[   49] = 'hb5048e03; 	    wvalid_rom[   49] = 0; 
    i_addr_rom[   50] = 'h000005bc; 	    d_addr_rom[   50] = 'h00000ce0; 	    wdata_rom[   50] = 'h53825215; 	    wvalid_rom[   50] = 1; 
    i_addr_rom[   51] = 'h00000374; 	    d_addr_rom[   51] = 'h000008b4; 	    wdata_rom[   51] = 'he1d50dc5; 	    wvalid_rom[   51] = 1; 
    i_addr_rom[   52] = 'h00000470; 	    d_addr_rom[   52] = 'h00000edc; 	    wdata_rom[   52] = 'h82f887b8; 	    wvalid_rom[   52] = 0; 
    i_addr_rom[   53] = 'h00000434; 	    d_addr_rom[   53] = 'h00000e4c; 	    wdata_rom[   53] = 'h3aa83c20; 	    wvalid_rom[   53] = 0; 
    i_addr_rom[   54] = 'h00000038; 	    d_addr_rom[   54] = 'h000009e0; 	    wdata_rom[   54] = 'h89868473; 	    wvalid_rom[   54] = 0; 
    i_addr_rom[   55] = 'h00000160; 	    d_addr_rom[   55] = 'h00000fd0; 	    wdata_rom[   55] = 'h89887f49; 	    wvalid_rom[   55] = 0; 
    i_addr_rom[   56] = 'h000006c8; 	    d_addr_rom[   56] = 'h00000c7c; 	    wdata_rom[   56] = 'h8ce85606; 	    wvalid_rom[   56] = 1; 
    i_addr_rom[   57] = 'h00000634; 	    d_addr_rom[   57] = 'h00000f2c; 	    wdata_rom[   57] = 'h6ca78010; 	    wvalid_rom[   57] = 0; 
    i_addr_rom[   58] = 'h000006bc; 	    d_addr_rom[   58] = 'h00000f10; 	    wdata_rom[   58] = 'h392aa1b7; 	    wvalid_rom[   58] = 1; 
    i_addr_rom[   59] = 'h00000568; 	    d_addr_rom[   59] = 'h00000c5c; 	    wdata_rom[   59] = 'hf64e7d72; 	    wvalid_rom[   59] = 1; 
    i_addr_rom[   60] = 'h00000268; 	    d_addr_rom[   60] = 'h00000c24; 	    wdata_rom[   60] = 'h04643dbe; 	    wvalid_rom[   60] = 1; 
    i_addr_rom[   61] = 'h00000294; 	    d_addr_rom[   61] = 'h00000c44; 	    wdata_rom[   61] = 'hbcf9b4d4; 	    wvalid_rom[   61] = 1; 
    i_addr_rom[   62] = 'h00000534; 	    d_addr_rom[   62] = 'h00000d94; 	    wdata_rom[   62] = 'ha978666d; 	    wvalid_rom[   62] = 0; 
    i_addr_rom[   63] = 'h00000744; 	    d_addr_rom[   63] = 'h00000934; 	    wdata_rom[   63] = 'h73cfa332; 	    wvalid_rom[   63] = 0; 
    i_addr_rom[   64] = 'h00000080; 	    d_addr_rom[   64] = 'h00000ed0; 	    wdata_rom[   64] = 'h6762f153; 	    wvalid_rom[   64] = 1; 
    i_addr_rom[   65] = 'h00000498; 	    d_addr_rom[   65] = 'h00000b00; 	    wdata_rom[   65] = 'h9f1e9983; 	    wvalid_rom[   65] = 0; 
    i_addr_rom[   66] = 'h000002cc; 	    d_addr_rom[   66] = 'h00000d6c; 	    wdata_rom[   66] = 'h5b3c9988; 	    wvalid_rom[   66] = 1; 
    i_addr_rom[   67] = 'h00000524; 	    d_addr_rom[   67] = 'h000009cc; 	    wdata_rom[   67] = 'h5bbfeb71; 	    wvalid_rom[   67] = 1; 
    i_addr_rom[   68] = 'h000006c0; 	    d_addr_rom[   68] = 'h00000a34; 	    wdata_rom[   68] = 'h77ec4a66; 	    wvalid_rom[   68] = 0; 
    i_addr_rom[   69] = 'h00000048; 	    d_addr_rom[   69] = 'h00000c94; 	    wdata_rom[   69] = 'hdcf9d6e5; 	    wvalid_rom[   69] = 1; 
    i_addr_rom[   70] = 'h000005a0; 	    d_addr_rom[   70] = 'h00000dbc; 	    wdata_rom[   70] = 'h506baa55; 	    wvalid_rom[   70] = 0; 
    i_addr_rom[   71] = 'h00000424; 	    d_addr_rom[   71] = 'h00000f78; 	    wdata_rom[   71] = 'h8a340fcc; 	    wvalid_rom[   71] = 0; 
    i_addr_rom[   72] = 'h00000050; 	    d_addr_rom[   72] = 'h00000a64; 	    wdata_rom[   72] = 'h02f9c470; 	    wvalid_rom[   72] = 0; 
    i_addr_rom[   73] = 'h000002d0; 	    d_addr_rom[   73] = 'h000009dc; 	    wdata_rom[   73] = 'h57f323ab; 	    wvalid_rom[   73] = 0; 
    i_addr_rom[   74] = 'h00000408; 	    d_addr_rom[   74] = 'h00000c20; 	    wdata_rom[   74] = 'ha03f3473; 	    wvalid_rom[   74] = 0; 
    i_addr_rom[   75] = 'h000007d8; 	    d_addr_rom[   75] = 'h00000dac; 	    wdata_rom[   75] = 'h677f5738; 	    wvalid_rom[   75] = 1; 
    i_addr_rom[   76] = 'h000002c4; 	    d_addr_rom[   76] = 'h00000e48; 	    wdata_rom[   76] = 'hdc8699b8; 	    wvalid_rom[   76] = 0; 
    i_addr_rom[   77] = 'h0000017c; 	    d_addr_rom[   77] = 'h00000b9c; 	    wdata_rom[   77] = 'hefbd668d; 	    wvalid_rom[   77] = 1; 
    i_addr_rom[   78] = 'h000006ac; 	    d_addr_rom[   78] = 'h00000bd0; 	    wdata_rom[   78] = 'hbafb8322; 	    wvalid_rom[   78] = 0; 
    i_addr_rom[   79] = 'h000001fc; 	    d_addr_rom[   79] = 'h0000080c; 	    wdata_rom[   79] = 'he131139e; 	    wvalid_rom[   79] = 0; 
    i_addr_rom[   80] = 'h000005c0; 	    d_addr_rom[   80] = 'h00000d1c; 	    wdata_rom[   80] = 'h8bb06312; 	    wvalid_rom[   80] = 0; 
    i_addr_rom[   81] = 'h000002d0; 	    d_addr_rom[   81] = 'h00000d2c; 	    wdata_rom[   81] = 'h8d00808c; 	    wvalid_rom[   81] = 0; 
    i_addr_rom[   82] = 'h000003ac; 	    d_addr_rom[   82] = 'h00000890; 	    wdata_rom[   82] = 'h11105786; 	    wvalid_rom[   82] = 0; 
    i_addr_rom[   83] = 'h00000370; 	    d_addr_rom[   83] = 'h00000d88; 	    wdata_rom[   83] = 'hebe69da3; 	    wvalid_rom[   83] = 1; 
    i_addr_rom[   84] = 'h000003a8; 	    d_addr_rom[   84] = 'h00000e34; 	    wdata_rom[   84] = 'hd29de744; 	    wvalid_rom[   84] = 0; 
    i_addr_rom[   85] = 'h00000500; 	    d_addr_rom[   85] = 'h00000900; 	    wdata_rom[   85] = 'h5c5a1e24; 	    wvalid_rom[   85] = 1; 
    i_addr_rom[   86] = 'h000002d0; 	    d_addr_rom[   86] = 'h00000d00; 	    wdata_rom[   86] = 'h32f63092; 	    wvalid_rom[   86] = 1; 
    i_addr_rom[   87] = 'h000003a4; 	    d_addr_rom[   87] = 'h00000ff8; 	    wdata_rom[   87] = 'hec78fedb; 	    wvalid_rom[   87] = 1; 
    i_addr_rom[   88] = 'h00000300; 	    d_addr_rom[   88] = 'h00000d1c; 	    wdata_rom[   88] = 'h211c3d36; 	    wvalid_rom[   88] = 1; 
    i_addr_rom[   89] = 'h00000790; 	    d_addr_rom[   89] = 'h00000ed4; 	    wdata_rom[   89] = 'h4048879c; 	    wvalid_rom[   89] = 0; 
    i_addr_rom[   90] = 'h0000065c; 	    d_addr_rom[   90] = 'h00000b70; 	    wdata_rom[   90] = 'h8c95cc91; 	    wvalid_rom[   90] = 1; 
    i_addr_rom[   91] = 'h00000594; 	    d_addr_rom[   91] = 'h00000ed4; 	    wdata_rom[   91] = 'h795c3538; 	    wvalid_rom[   91] = 1; 
    i_addr_rom[   92] = 'h00000264; 	    d_addr_rom[   92] = 'h000009a8; 	    wdata_rom[   92] = 'hd79766c1; 	    wvalid_rom[   92] = 1; 
    i_addr_rom[   93] = 'h000002cc; 	    d_addr_rom[   93] = 'h0000082c; 	    wdata_rom[   93] = 'hd04d3c52; 	    wvalid_rom[   93] = 0; 
    i_addr_rom[   94] = 'h00000164; 	    d_addr_rom[   94] = 'h00000c40; 	    wdata_rom[   94] = 'habd1db13; 	    wvalid_rom[   94] = 1; 
    i_addr_rom[   95] = 'h00000688; 	    d_addr_rom[   95] = 'h00000e9c; 	    wdata_rom[   95] = 'hc07774e8; 	    wvalid_rom[   95] = 0; 
    i_addr_rom[   96] = 'h000003fc; 	    d_addr_rom[   96] = 'h00000cb0; 	    wdata_rom[   96] = 'h91016ef2; 	    wvalid_rom[   96] = 1; 
    i_addr_rom[   97] = 'h0000055c; 	    d_addr_rom[   97] = 'h00000984; 	    wdata_rom[   97] = 'hc29daccd; 	    wvalid_rom[   97] = 1; 
    i_addr_rom[   98] = 'h00000698; 	    d_addr_rom[   98] = 'h00000b9c; 	    wdata_rom[   98] = 'h47ace802; 	    wvalid_rom[   98] = 1; 
    i_addr_rom[   99] = 'h00000220; 	    d_addr_rom[   99] = 'h00000f98; 	    wdata_rom[   99] = 'h2a57abb5; 	    wvalid_rom[   99] = 1; 
    i_addr_rom[  100] = 'h00000528; 	    d_addr_rom[  100] = 'h00000fd4; 	    wdata_rom[  100] = 'h0a822345; 	    wvalid_rom[  100] = 0; 
    i_addr_rom[  101] = 'h00000000; 	    d_addr_rom[  101] = 'h00000c44; 	    wdata_rom[  101] = 'h585915be; 	    wvalid_rom[  101] = 0; 
    i_addr_rom[  102] = 'h000003c8; 	    d_addr_rom[  102] = 'h00000ac8; 	    wdata_rom[  102] = 'h218dfe8d; 	    wvalid_rom[  102] = 0; 
    i_addr_rom[  103] = 'h000000f0; 	    d_addr_rom[  103] = 'h00000b5c; 	    wdata_rom[  103] = 'h5ceee06b; 	    wvalid_rom[  103] = 0; 
    i_addr_rom[  104] = 'h00000638; 	    d_addr_rom[  104] = 'h00000d54; 	    wdata_rom[  104] = 'h10ed02a7; 	    wvalid_rom[  104] = 0; 
    i_addr_rom[  105] = 'h00000554; 	    d_addr_rom[  105] = 'h00000fe4; 	    wdata_rom[  105] = 'h9fc5204b; 	    wvalid_rom[  105] = 1; 
    i_addr_rom[  106] = 'h00000690; 	    d_addr_rom[  106] = 'h00000e60; 	    wdata_rom[  106] = 'h0f35475b; 	    wvalid_rom[  106] = 1; 
    i_addr_rom[  107] = 'h0000057c; 	    d_addr_rom[  107] = 'h0000092c; 	    wdata_rom[  107] = 'h649679ba; 	    wvalid_rom[  107] = 1; 
    i_addr_rom[  108] = 'h000007d0; 	    d_addr_rom[  108] = 'h00000958; 	    wdata_rom[  108] = 'h1f99c3e1; 	    wvalid_rom[  108] = 1; 
    i_addr_rom[  109] = 'h0000055c; 	    d_addr_rom[  109] = 'h00000fa4; 	    wdata_rom[  109] = 'hcda7806f; 	    wvalid_rom[  109] = 1; 
    i_addr_rom[  110] = 'h0000012c; 	    d_addr_rom[  110] = 'h00000fc0; 	    wdata_rom[  110] = 'h3d367161; 	    wvalid_rom[  110] = 1; 
    i_addr_rom[  111] = 'h00000258; 	    d_addr_rom[  111] = 'h00000b2c; 	    wdata_rom[  111] = 'h84df8e45; 	    wvalid_rom[  111] = 0; 
    i_addr_rom[  112] = 'h0000068c; 	    d_addr_rom[  112] = 'h00000f20; 	    wdata_rom[  112] = 'h7fb3a30d; 	    wvalid_rom[  112] = 0; 
    i_addr_rom[  113] = 'h000001fc; 	    d_addr_rom[  113] = 'h00000eb4; 	    wdata_rom[  113] = 'hb1f3e1e5; 	    wvalid_rom[  113] = 0; 
    i_addr_rom[  114] = 'h00000140; 	    d_addr_rom[  114] = 'h000009e4; 	    wdata_rom[  114] = 'he395ceca; 	    wvalid_rom[  114] = 0; 
    i_addr_rom[  115] = 'h00000590; 	    d_addr_rom[  115] = 'h00000f3c; 	    wdata_rom[  115] = 'he5cb21d0; 	    wvalid_rom[  115] = 0; 
    i_addr_rom[  116] = 'h0000040c; 	    d_addr_rom[  116] = 'h0000088c; 	    wdata_rom[  116] = 'hbe90d535; 	    wvalid_rom[  116] = 0; 
    i_addr_rom[  117] = 'h000005a4; 	    d_addr_rom[  117] = 'h00000ab0; 	    wdata_rom[  117] = 'hba66255f; 	    wvalid_rom[  117] = 1; 
    i_addr_rom[  118] = 'h000003e8; 	    d_addr_rom[  118] = 'h00000d38; 	    wdata_rom[  118] = 'h7537a3b2; 	    wvalid_rom[  118] = 0; 
    i_addr_rom[  119] = 'h00000410; 	    d_addr_rom[  119] = 'h00000dac; 	    wdata_rom[  119] = 'h5407f98b; 	    wvalid_rom[  119] = 0; 
    i_addr_rom[  120] = 'h0000008c; 	    d_addr_rom[  120] = 'h00000ee4; 	    wdata_rom[  120] = 'h50142dcc; 	    wvalid_rom[  120] = 0; 
    i_addr_rom[  121] = 'h0000031c; 	    d_addr_rom[  121] = 'h00000f98; 	    wdata_rom[  121] = 'h390c7ff2; 	    wvalid_rom[  121] = 0; 
    i_addr_rom[  122] = 'h000004e4; 	    d_addr_rom[  122] = 'h000009bc; 	    wdata_rom[  122] = 'h1dd25d45; 	    wvalid_rom[  122] = 0; 
    i_addr_rom[  123] = 'h000001d8; 	    d_addr_rom[  123] = 'h000009d4; 	    wdata_rom[  123] = 'h9e99f3f3; 	    wvalid_rom[  123] = 0; 
    i_addr_rom[  124] = 'h00000538; 	    d_addr_rom[  124] = 'h00000b70; 	    wdata_rom[  124] = 'h74e43485; 	    wvalid_rom[  124] = 1; 
    i_addr_rom[  125] = 'h0000006c; 	    d_addr_rom[  125] = 'h00000eec; 	    wdata_rom[  125] = 'h55e9ab61; 	    wvalid_rom[  125] = 1; 
    i_addr_rom[  126] = 'h00000488; 	    d_addr_rom[  126] = 'h00000cd8; 	    wdata_rom[  126] = 'h06ee75e3; 	    wvalid_rom[  126] = 1; 
    i_addr_rom[  127] = 'h000001cc; 	    d_addr_rom[  127] = 'h00000b74; 	    wdata_rom[  127] = 'h44a66839; 	    wvalid_rom[  127] = 1; 
    i_addr_rom[  128] = 'h0000015c; 	    d_addr_rom[  128] = 'h00000ea4; 	    wdata_rom[  128] = 'h1f076333; 	    wvalid_rom[  128] = 1; 
    i_addr_rom[  129] = 'h000006e4; 	    d_addr_rom[  129] = 'h000008c4; 	    wdata_rom[  129] = 'h59a8ff6c; 	    wvalid_rom[  129] = 1; 
    i_addr_rom[  130] = 'h000003b0; 	    d_addr_rom[  130] = 'h00000fac; 	    wdata_rom[  130] = 'ha9fe429e; 	    wvalid_rom[  130] = 0; 
    i_addr_rom[  131] = 'h00000774; 	    d_addr_rom[  131] = 'h00000cec; 	    wdata_rom[  131] = 'h880e2269; 	    wvalid_rom[  131] = 1; 
    i_addr_rom[  132] = 'h0000002c; 	    d_addr_rom[  132] = 'h00000c74; 	    wdata_rom[  132] = 'hb2aa5851; 	    wvalid_rom[  132] = 0; 
    i_addr_rom[  133] = 'h00000488; 	    d_addr_rom[  133] = 'h00000f18; 	    wdata_rom[  133] = 'h31ecc96b; 	    wvalid_rom[  133] = 1; 
    i_addr_rom[  134] = 'h0000027c; 	    d_addr_rom[  134] = 'h00000ed8; 	    wdata_rom[  134] = 'h0ae71fe2; 	    wvalid_rom[  134] = 1; 
    i_addr_rom[  135] = 'h00000390; 	    d_addr_rom[  135] = 'h00000d68; 	    wdata_rom[  135] = 'he50a491f; 	    wvalid_rom[  135] = 0; 
    i_addr_rom[  136] = 'h0000067c; 	    d_addr_rom[  136] = 'h00000b18; 	    wdata_rom[  136] = 'h5b52bed3; 	    wvalid_rom[  136] = 0; 
    i_addr_rom[  137] = 'h0000026c; 	    d_addr_rom[  137] = 'h00000ef4; 	    wdata_rom[  137] = 'haed7b3fb; 	    wvalid_rom[  137] = 1; 
    i_addr_rom[  138] = 'h00000168; 	    d_addr_rom[  138] = 'h00000870; 	    wdata_rom[  138] = 'haafa909b; 	    wvalid_rom[  138] = 0; 
    i_addr_rom[  139] = 'h0000066c; 	    d_addr_rom[  139] = 'h00000b48; 	    wdata_rom[  139] = 'h41745b6b; 	    wvalid_rom[  139] = 0; 
    i_addr_rom[  140] = 'h000003b4; 	    d_addr_rom[  140] = 'h00000958; 	    wdata_rom[  140] = 'hc65bb258; 	    wvalid_rom[  140] = 1; 
    i_addr_rom[  141] = 'h000002ac; 	    d_addr_rom[  141] = 'h00000ce4; 	    wdata_rom[  141] = 'hedb7db79; 	    wvalid_rom[  141] = 1; 
    i_addr_rom[  142] = 'h000003dc; 	    d_addr_rom[  142] = 'h00000918; 	    wdata_rom[  142] = 'he4db56dc; 	    wvalid_rom[  142] = 1; 
    i_addr_rom[  143] = 'h00000754; 	    d_addr_rom[  143] = 'h00000cac; 	    wdata_rom[  143] = 'h21cec50d; 	    wvalid_rom[  143] = 1; 
    i_addr_rom[  144] = 'h000004e0; 	    d_addr_rom[  144] = 'h00000ec0; 	    wdata_rom[  144] = 'h4fbba5fe; 	    wvalid_rom[  144] = 0; 
    i_addr_rom[  145] = 'h000007c8; 	    d_addr_rom[  145] = 'h0000080c; 	    wdata_rom[  145] = 'hef6c0d43; 	    wvalid_rom[  145] = 0; 
    i_addr_rom[  146] = 'h00000798; 	    d_addr_rom[  146] = 'h00000bc0; 	    wdata_rom[  146] = 'h20c59047; 	    wvalid_rom[  146] = 0; 
    i_addr_rom[  147] = 'h00000530; 	    d_addr_rom[  147] = 'h000008b0; 	    wdata_rom[  147] = 'h6d52ef58; 	    wvalid_rom[  147] = 1; 
    i_addr_rom[  148] = 'h00000614; 	    d_addr_rom[  148] = 'h00000c50; 	    wdata_rom[  148] = 'he1f61c9d; 	    wvalid_rom[  148] = 1; 
    i_addr_rom[  149] = 'h000000f0; 	    d_addr_rom[  149] = 'h00000d60; 	    wdata_rom[  149] = 'hf5eb38e9; 	    wvalid_rom[  149] = 1; 
    i_addr_rom[  150] = 'h000007c8; 	    d_addr_rom[  150] = 'h00000fb0; 	    wdata_rom[  150] = 'he3eab3e1; 	    wvalid_rom[  150] = 0; 
    i_addr_rom[  151] = 'h00000294; 	    d_addr_rom[  151] = 'h00000b48; 	    wdata_rom[  151] = 'he1e26668; 	    wvalid_rom[  151] = 1; 
    i_addr_rom[  152] = 'h00000180; 	    d_addr_rom[  152] = 'h00000ff0; 	    wdata_rom[  152] = 'h89ca9bf4; 	    wvalid_rom[  152] = 0; 
    i_addr_rom[  153] = 'h000006a4; 	    d_addr_rom[  153] = 'h00000810; 	    wdata_rom[  153] = 'hb1dfdd87; 	    wvalid_rom[  153] = 1; 
    i_addr_rom[  154] = 'h00000750; 	    d_addr_rom[  154] = 'h00000fd4; 	    wdata_rom[  154] = 'h9fa8b417; 	    wvalid_rom[  154] = 1; 
    i_addr_rom[  155] = 'h00000010; 	    d_addr_rom[  155] = 'h00000aa4; 	    wdata_rom[  155] = 'hec9c72cb; 	    wvalid_rom[  155] = 0; 
    i_addr_rom[  156] = 'h000002a8; 	    d_addr_rom[  156] = 'h00000acc; 	    wdata_rom[  156] = 'h7724aff5; 	    wvalid_rom[  156] = 1; 
    i_addr_rom[  157] = 'h00000574; 	    d_addr_rom[  157] = 'h00000970; 	    wdata_rom[  157] = 'hd132e7bb; 	    wvalid_rom[  157] = 1; 
    i_addr_rom[  158] = 'h00000610; 	    d_addr_rom[  158] = 'h00000d04; 	    wdata_rom[  158] = 'h628c539f; 	    wvalid_rom[  158] = 0; 
    i_addr_rom[  159] = 'h00000308; 	    d_addr_rom[  159] = 'h00000bd0; 	    wdata_rom[  159] = 'h54dd8c4e; 	    wvalid_rom[  159] = 0; 
    i_addr_rom[  160] = 'h0000075c; 	    d_addr_rom[  160] = 'h00000c80; 	    wdata_rom[  160] = 'haf45c266; 	    wvalid_rom[  160] = 0; 
    i_addr_rom[  161] = 'h000001cc; 	    d_addr_rom[  161] = 'h00000da0; 	    wdata_rom[  161] = 'h81bb4f51; 	    wvalid_rom[  161] = 0; 
    i_addr_rom[  162] = 'h00000120; 	    d_addr_rom[  162] = 'h00000f88; 	    wdata_rom[  162] = 'h7619d9a9; 	    wvalid_rom[  162] = 1; 
    i_addr_rom[  163] = 'h000004f0; 	    d_addr_rom[  163] = 'h00000f60; 	    wdata_rom[  163] = 'habf1f234; 	    wvalid_rom[  163] = 0; 
    i_addr_rom[  164] = 'h00000044; 	    d_addr_rom[  164] = 'h00000aec; 	    wdata_rom[  164] = 'hcb3d120a; 	    wvalid_rom[  164] = 1; 
    i_addr_rom[  165] = 'h00000354; 	    d_addr_rom[  165] = 'h0000097c; 	    wdata_rom[  165] = 'heef6283c; 	    wvalid_rom[  165] = 1; 
    i_addr_rom[  166] = 'h0000043c; 	    d_addr_rom[  166] = 'h0000083c; 	    wdata_rom[  166] = 'hbd9391be; 	    wvalid_rom[  166] = 0; 
    i_addr_rom[  167] = 'h0000018c; 	    d_addr_rom[  167] = 'h00000814; 	    wdata_rom[  167] = 'h4aaf2bc3; 	    wvalid_rom[  167] = 1; 
    i_addr_rom[  168] = 'h0000068c; 	    d_addr_rom[  168] = 'h00000aa8; 	    wdata_rom[  168] = 'ha2cddaed; 	    wvalid_rom[  168] = 0; 
    i_addr_rom[  169] = 'h0000005c; 	    d_addr_rom[  169] = 'h00000bec; 	    wdata_rom[  169] = 'h02b910c9; 	    wvalid_rom[  169] = 1; 
    i_addr_rom[  170] = 'h000007a4; 	    d_addr_rom[  170] = 'h00000c78; 	    wdata_rom[  170] = 'h1a3b8ae6; 	    wvalid_rom[  170] = 1; 
    i_addr_rom[  171] = 'h0000068c; 	    d_addr_rom[  171] = 'h00000a90; 	    wdata_rom[  171] = 'h708019a9; 	    wvalid_rom[  171] = 0; 
    i_addr_rom[  172] = 'h00000280; 	    d_addr_rom[  172] = 'h000009b8; 	    wdata_rom[  172] = 'h433defb5; 	    wvalid_rom[  172] = 1; 
    i_addr_rom[  173] = 'h000002b8; 	    d_addr_rom[  173] = 'h00000dfc; 	    wdata_rom[  173] = 'h049e3fd7; 	    wvalid_rom[  173] = 1; 
    i_addr_rom[  174] = 'h00000230; 	    d_addr_rom[  174] = 'h00000fb0; 	    wdata_rom[  174] = 'h02f5adce; 	    wvalid_rom[  174] = 0; 
    i_addr_rom[  175] = 'h00000310; 	    d_addr_rom[  175] = 'h00000e1c; 	    wdata_rom[  175] = 'he27069a7; 	    wvalid_rom[  175] = 1; 
    i_addr_rom[  176] = 'h000007a8; 	    d_addr_rom[  176] = 'h00000a20; 	    wdata_rom[  176] = 'h4b9fa00f; 	    wvalid_rom[  176] = 1; 
    i_addr_rom[  177] = 'h000006ec; 	    d_addr_rom[  177] = 'h00000a34; 	    wdata_rom[  177] = 'h05600812; 	    wvalid_rom[  177] = 1; 
    i_addr_rom[  178] = 'h000000dc; 	    d_addr_rom[  178] = 'h00000a18; 	    wdata_rom[  178] = 'h81fcd450; 	    wvalid_rom[  178] = 1; 
    i_addr_rom[  179] = 'h00000568; 	    d_addr_rom[  179] = 'h00000d1c; 	    wdata_rom[  179] = 'h8fb3f291; 	    wvalid_rom[  179] = 0; 
    i_addr_rom[  180] = 'h00000328; 	    d_addr_rom[  180] = 'h00000ca8; 	    wdata_rom[  180] = 'hedca4df1; 	    wvalid_rom[  180] = 0; 
    i_addr_rom[  181] = 'h00000080; 	    d_addr_rom[  181] = 'h00000990; 	    wdata_rom[  181] = 'hf272cb6d; 	    wvalid_rom[  181] = 1; 
    i_addr_rom[  182] = 'h00000364; 	    d_addr_rom[  182] = 'h00000bb4; 	    wdata_rom[  182] = 'h9d6bf2e4; 	    wvalid_rom[  182] = 0; 
    i_addr_rom[  183] = 'h000004d8; 	    d_addr_rom[  183] = 'h00000970; 	    wdata_rom[  183] = 'h8ec460af; 	    wvalid_rom[  183] = 0; 
    i_addr_rom[  184] = 'h0000036c; 	    d_addr_rom[  184] = 'h00000d0c; 	    wdata_rom[  184] = 'h9a1e1ab7; 	    wvalid_rom[  184] = 1; 
    i_addr_rom[  185] = 'h0000038c; 	    d_addr_rom[  185] = 'h000009a4; 	    wdata_rom[  185] = 'h4074788a; 	    wvalid_rom[  185] = 0; 
    i_addr_rom[  186] = 'h000000fc; 	    d_addr_rom[  186] = 'h00000e80; 	    wdata_rom[  186] = 'hc561154f; 	    wvalid_rom[  186] = 0; 
    i_addr_rom[  187] = 'h000007cc; 	    d_addr_rom[  187] = 'h00000c2c; 	    wdata_rom[  187] = 'h10c02679; 	    wvalid_rom[  187] = 1; 
    i_addr_rom[  188] = 'h000003fc; 	    d_addr_rom[  188] = 'h000009b8; 	    wdata_rom[  188] = 'h8ee2523c; 	    wvalid_rom[  188] = 0; 
    i_addr_rom[  189] = 'h000003b0; 	    d_addr_rom[  189] = 'h00000bc4; 	    wdata_rom[  189] = 'h9d921cdc; 	    wvalid_rom[  189] = 0; 
    i_addr_rom[  190] = 'h00000638; 	    d_addr_rom[  190] = 'h00000c1c; 	    wdata_rom[  190] = 'hf1fbd347; 	    wvalid_rom[  190] = 0; 
    i_addr_rom[  191] = 'h000000b4; 	    d_addr_rom[  191] = 'h00000934; 	    wdata_rom[  191] = 'hc99dc9aa; 	    wvalid_rom[  191] = 0; 
    i_addr_rom[  192] = 'h00000720; 	    d_addr_rom[  192] = 'h00000d54; 	    wdata_rom[  192] = 'hec16b630; 	    wvalid_rom[  192] = 0; 
    i_addr_rom[  193] = 'h0000021c; 	    d_addr_rom[  193] = 'h00000b0c; 	    wdata_rom[  193] = 'h1657b4af; 	    wvalid_rom[  193] = 1; 
    i_addr_rom[  194] = 'h00000454; 	    d_addr_rom[  194] = 'h00000b0c; 	    wdata_rom[  194] = 'hcf550517; 	    wvalid_rom[  194] = 1; 
    i_addr_rom[  195] = 'h0000017c; 	    d_addr_rom[  195] = 'h00000ab4; 	    wdata_rom[  195] = 'h12afc44a; 	    wvalid_rom[  195] = 0; 
    i_addr_rom[  196] = 'h000003a8; 	    d_addr_rom[  196] = 'h00000d64; 	    wdata_rom[  196] = 'h80851384; 	    wvalid_rom[  196] = 1; 
    i_addr_rom[  197] = 'h000006ec; 	    d_addr_rom[  197] = 'h00000ee8; 	    wdata_rom[  197] = 'h690e0c39; 	    wvalid_rom[  197] = 0; 
    i_addr_rom[  198] = 'h00000484; 	    d_addr_rom[  198] = 'h00000aa4; 	    wdata_rom[  198] = 'h0386f463; 	    wvalid_rom[  198] = 1; 
    i_addr_rom[  199] = 'h00000798; 	    d_addr_rom[  199] = 'h00000ea8; 	    wdata_rom[  199] = 'h816132aa; 	    wvalid_rom[  199] = 0; 
    i_addr_rom[  200] = 'h00000608; 	    d_addr_rom[  200] = 'h00000914; 	    wdata_rom[  200] = 'hd8dc6984; 	    wvalid_rom[  200] = 1; 
    i_addr_rom[  201] = 'h00000098; 	    d_addr_rom[  201] = 'h00000f24; 	    wdata_rom[  201] = 'hcb30120e; 	    wvalid_rom[  201] = 1; 
    i_addr_rom[  202] = 'h0000052c; 	    d_addr_rom[  202] = 'h00000e1c; 	    wdata_rom[  202] = 'h53a30946; 	    wvalid_rom[  202] = 0; 
    i_addr_rom[  203] = 'h00000524; 	    d_addr_rom[  203] = 'h00000c10; 	    wdata_rom[  203] = 'h5233804c; 	    wvalid_rom[  203] = 0; 
    i_addr_rom[  204] = 'h00000414; 	    d_addr_rom[  204] = 'h00000b48; 	    wdata_rom[  204] = 'h3e68c860; 	    wvalid_rom[  204] = 1; 
    i_addr_rom[  205] = 'h000003fc; 	    d_addr_rom[  205] = 'h00000c9c; 	    wdata_rom[  205] = 'hf86aecce; 	    wvalid_rom[  205] = 0; 
    i_addr_rom[  206] = 'h00000320; 	    d_addr_rom[  206] = 'h00000d78; 	    wdata_rom[  206] = 'h616f7e76; 	    wvalid_rom[  206] = 0; 
    i_addr_rom[  207] = 'h000005b0; 	    d_addr_rom[  207] = 'h00000b2c; 	    wdata_rom[  207] = 'h4b6e80fb; 	    wvalid_rom[  207] = 1; 
    i_addr_rom[  208] = 'h000001cc; 	    d_addr_rom[  208] = 'h00000ddc; 	    wdata_rom[  208] = 'h2d838389; 	    wvalid_rom[  208] = 0; 
    i_addr_rom[  209] = 'h00000498; 	    d_addr_rom[  209] = 'h00000e78; 	    wdata_rom[  209] = 'h9f7fea57; 	    wvalid_rom[  209] = 1; 
    i_addr_rom[  210] = 'h00000788; 	    d_addr_rom[  210] = 'h00000d84; 	    wdata_rom[  210] = 'h371ab284; 	    wvalid_rom[  210] = 1; 
    i_addr_rom[  211] = 'h000000f4; 	    d_addr_rom[  211] = 'h000008c4; 	    wdata_rom[  211] = 'hc3e30f5b; 	    wvalid_rom[  211] = 1; 
    i_addr_rom[  212] = 'h000005f8; 	    d_addr_rom[  212] = 'h000009c8; 	    wdata_rom[  212] = 'he2677277; 	    wvalid_rom[  212] = 0; 
    i_addr_rom[  213] = 'h000005d8; 	    d_addr_rom[  213] = 'h00000df4; 	    wdata_rom[  213] = 'h823c59f6; 	    wvalid_rom[  213] = 0; 
    i_addr_rom[  214] = 'h000006cc; 	    d_addr_rom[  214] = 'h00000fb4; 	    wdata_rom[  214] = 'h9c6212bd; 	    wvalid_rom[  214] = 0; 
    i_addr_rom[  215] = 'h00000458; 	    d_addr_rom[  215] = 'h00000e74; 	    wdata_rom[  215] = 'hc3c869fa; 	    wvalid_rom[  215] = 0; 
    i_addr_rom[  216] = 'h000005c8; 	    d_addr_rom[  216] = 'h00000eb4; 	    wdata_rom[  216] = 'hf5272cbf; 	    wvalid_rom[  216] = 1; 
    i_addr_rom[  217] = 'h00000248; 	    d_addr_rom[  217] = 'h00000aa0; 	    wdata_rom[  217] = 'hfe29a2e6; 	    wvalid_rom[  217] = 0; 
    i_addr_rom[  218] = 'h00000598; 	    d_addr_rom[  218] = 'h00000a40; 	    wdata_rom[  218] = 'h74f5f8f0; 	    wvalid_rom[  218] = 0; 
    i_addr_rom[  219] = 'h000001b8; 	    d_addr_rom[  219] = 'h00000fb0; 	    wdata_rom[  219] = 'hc47f475f; 	    wvalid_rom[  219] = 0; 
    i_addr_rom[  220] = 'h000005f8; 	    d_addr_rom[  220] = 'h000009c0; 	    wdata_rom[  220] = 'h1eb5bde1; 	    wvalid_rom[  220] = 0; 
    i_addr_rom[  221] = 'h000000bc; 	    d_addr_rom[  221] = 'h00000d20; 	    wdata_rom[  221] = 'h5b90d8a9; 	    wvalid_rom[  221] = 1; 
    i_addr_rom[  222] = 'h000005d8; 	    d_addr_rom[  222] = 'h00000f20; 	    wdata_rom[  222] = 'h08c4d7fc; 	    wvalid_rom[  222] = 0; 
    i_addr_rom[  223] = 'h00000080; 	    d_addr_rom[  223] = 'h00000bb4; 	    wdata_rom[  223] = 'h0238be6c; 	    wvalid_rom[  223] = 0; 
    i_addr_rom[  224] = 'h00000298; 	    d_addr_rom[  224] = 'h000008fc; 	    wdata_rom[  224] = 'h1fde48f6; 	    wvalid_rom[  224] = 0; 
    i_addr_rom[  225] = 'h0000070c; 	    d_addr_rom[  225] = 'h000008e8; 	    wdata_rom[  225] = 'hae78e1ce; 	    wvalid_rom[  225] = 0; 
    i_addr_rom[  226] = 'h000001b4; 	    d_addr_rom[  226] = 'h00000a60; 	    wdata_rom[  226] = 'hb57e362a; 	    wvalid_rom[  226] = 1; 
    i_addr_rom[  227] = 'h000005f8; 	    d_addr_rom[  227] = 'h00000dcc; 	    wdata_rom[  227] = 'ha6827dd6; 	    wvalid_rom[  227] = 1; 
    i_addr_rom[  228] = 'h00000328; 	    d_addr_rom[  228] = 'h00000db4; 	    wdata_rom[  228] = 'ha5112ecc; 	    wvalid_rom[  228] = 1; 
    i_addr_rom[  229] = 'h000005e8; 	    d_addr_rom[  229] = 'h00000fe0; 	    wdata_rom[  229] = 'haeb5305e; 	    wvalid_rom[  229] = 0; 
    i_addr_rom[  230] = 'h000004fc; 	    d_addr_rom[  230] = 'h00000f0c; 	    wdata_rom[  230] = 'he8a531ab; 	    wvalid_rom[  230] = 1; 
    i_addr_rom[  231] = 'h000000a8; 	    d_addr_rom[  231] = 'h000009dc; 	    wdata_rom[  231] = 'hff8d6edf; 	    wvalid_rom[  231] = 1; 
    i_addr_rom[  232] = 'h000000b0; 	    d_addr_rom[  232] = 'h00000924; 	    wdata_rom[  232] = 'h05fb3028; 	    wvalid_rom[  232] = 1; 
    i_addr_rom[  233] = 'h000005b8; 	    d_addr_rom[  233] = 'h00000bc8; 	    wdata_rom[  233] = 'hc83a8ab6; 	    wvalid_rom[  233] = 0; 
    i_addr_rom[  234] = 'h000007cc; 	    d_addr_rom[  234] = 'h00000b74; 	    wdata_rom[  234] = 'h92839366; 	    wvalid_rom[  234] = 1; 
    i_addr_rom[  235] = 'h00000268; 	    d_addr_rom[  235] = 'h00000b6c; 	    wdata_rom[  235] = 'haa169388; 	    wvalid_rom[  235] = 1; 
    i_addr_rom[  236] = 'h000000e8; 	    d_addr_rom[  236] = 'h00000b0c; 	    wdata_rom[  236] = 'h8ed6c144; 	    wvalid_rom[  236] = 1; 
    i_addr_rom[  237] = 'h000004d8; 	    d_addr_rom[  237] = 'h000008b0; 	    wdata_rom[  237] = 'hd17c2b5a; 	    wvalid_rom[  237] = 1; 
    i_addr_rom[  238] = 'h00000560; 	    d_addr_rom[  238] = 'h0000097c; 	    wdata_rom[  238] = 'h451db60d; 	    wvalid_rom[  238] = 0; 
    i_addr_rom[  239] = 'h00000310; 	    d_addr_rom[  239] = 'h000008ac; 	    wdata_rom[  239] = 'h8e2e7384; 	    wvalid_rom[  239] = 0; 
    i_addr_rom[  240] = 'h00000288; 	    d_addr_rom[  240] = 'h0000080c; 	    wdata_rom[  240] = 'h77482af6; 	    wvalid_rom[  240] = 1; 
    i_addr_rom[  241] = 'h00000350; 	    d_addr_rom[  241] = 'h00000d00; 	    wdata_rom[  241] = 'hdfc87209; 	    wvalid_rom[  241] = 0; 
    i_addr_rom[  242] = 'h00000348; 	    d_addr_rom[  242] = 'h00000ae4; 	    wdata_rom[  242] = 'h82d222b3; 	    wvalid_rom[  242] = 1; 
    i_addr_rom[  243] = 'h00000550; 	    d_addr_rom[  243] = 'h00000d6c; 	    wdata_rom[  243] = 'he3ffb632; 	    wvalid_rom[  243] = 1; 
    i_addr_rom[  244] = 'h000006a8; 	    d_addr_rom[  244] = 'h00000914; 	    wdata_rom[  244] = 'h37c7da1e; 	    wvalid_rom[  244] = 1; 
    i_addr_rom[  245] = 'h00000500; 	    d_addr_rom[  245] = 'h00000f38; 	    wdata_rom[  245] = 'h9b5ae3d7; 	    wvalid_rom[  245] = 0; 
    i_addr_rom[  246] = 'h00000128; 	    d_addr_rom[  246] = 'h000008ec; 	    wdata_rom[  246] = 'heb488c96; 	    wvalid_rom[  246] = 1; 
    i_addr_rom[  247] = 'h000004fc; 	    d_addr_rom[  247] = 'h00000a20; 	    wdata_rom[  247] = 'h541a37a3; 	    wvalid_rom[  247] = 0; 
    i_addr_rom[  248] = 'h00000110; 	    d_addr_rom[  248] = 'h00000bcc; 	    wdata_rom[  248] = 'h2e883bc5; 	    wvalid_rom[  248] = 1; 
    i_addr_rom[  249] = 'h00000648; 	    d_addr_rom[  249] = 'h00000e30; 	    wdata_rom[  249] = 'h8fe2c67d; 	    wvalid_rom[  249] = 1; 
    i_addr_rom[  250] = 'h000002d0; 	    d_addr_rom[  250] = 'h00000de0; 	    wdata_rom[  250] = 'hf8dc2f83; 	    wvalid_rom[  250] = 0; 
    i_addr_rom[  251] = 'h000007ec; 	    d_addr_rom[  251] = 'h00000aa4; 	    wdata_rom[  251] = 'hd4cffbf9; 	    wvalid_rom[  251] = 1; 
    i_addr_rom[  252] = 'h00000678; 	    d_addr_rom[  252] = 'h0000097c; 	    wdata_rom[  252] = 'hcbc49136; 	    wvalid_rom[  252] = 1; 
    i_addr_rom[  253] = 'h000005b4; 	    d_addr_rom[  253] = 'h00000bf0; 	    wdata_rom[  253] = 'hea87f38f; 	    wvalid_rom[  253] = 1; 
    i_addr_rom[  254] = 'h000006b0; 	    d_addr_rom[  254] = 'h00000a44; 	    wdata_rom[  254] = 'h22f9f4a2; 	    wvalid_rom[  254] = 0; 
    i_addr_rom[  255] = 'h000003cc; 	    d_addr_rom[  255] = 'h00000db8; 	    wdata_rom[  255] = 'hf6f7fd01; 	    wvalid_rom[  255] = 0; 
    i_addr_rom[  256] = 'h00000180; 	    d_addr_rom[  256] = 'h00000ffc; 	    wdata_rom[  256] = 'he6b84af2; 	    wvalid_rom[  256] = 0; 
    i_addr_rom[  257] = 'h0000025c; 	    d_addr_rom[  257] = 'h00000ea0; 	    wdata_rom[  257] = 'hbd4fc407; 	    wvalid_rom[  257] = 1; 
    i_addr_rom[  258] = 'h00000580; 	    d_addr_rom[  258] = 'h00000cc8; 	    wdata_rom[  258] = 'h81d20e16; 	    wvalid_rom[  258] = 0; 
    i_addr_rom[  259] = 'h00000070; 	    d_addr_rom[  259] = 'h00000dec; 	    wdata_rom[  259] = 'h2ac199df; 	    wvalid_rom[  259] = 0; 
    i_addr_rom[  260] = 'h00000504; 	    d_addr_rom[  260] = 'h00000e6c; 	    wdata_rom[  260] = 'hb33f0cf2; 	    wvalid_rom[  260] = 0; 
    i_addr_rom[  261] = 'h00000350; 	    d_addr_rom[  261] = 'h00000e9c; 	    wdata_rom[  261] = 'h5f2f5e69; 	    wvalid_rom[  261] = 1; 
    i_addr_rom[  262] = 'h00000318; 	    d_addr_rom[  262] = 'h00000d54; 	    wdata_rom[  262] = 'hcae66eb7; 	    wvalid_rom[  262] = 1; 
    i_addr_rom[  263] = 'h00000770; 	    d_addr_rom[  263] = 'h00000c88; 	    wdata_rom[  263] = 'h928e3138; 	    wvalid_rom[  263] = 1; 
    i_addr_rom[  264] = 'h0000079c; 	    d_addr_rom[  264] = 'h00000928; 	    wdata_rom[  264] = 'hbe83cd02; 	    wvalid_rom[  264] = 0; 
    i_addr_rom[  265] = 'h000001c0; 	    d_addr_rom[  265] = 'h00000bb8; 	    wdata_rom[  265] = 'hab8e4dfa; 	    wvalid_rom[  265] = 1; 
    i_addr_rom[  266] = 'h00000118; 	    d_addr_rom[  266] = 'h00000aa0; 	    wdata_rom[  266] = 'h9dac9b9c; 	    wvalid_rom[  266] = 0; 
    i_addr_rom[  267] = 'h0000031c; 	    d_addr_rom[  267] = 'h00000aa8; 	    wdata_rom[  267] = 'h0727b204; 	    wvalid_rom[  267] = 0; 
    i_addr_rom[  268] = 'h00000190; 	    d_addr_rom[  268] = 'h00000a68; 	    wdata_rom[  268] = 'h0b40f5ba; 	    wvalid_rom[  268] = 1; 
    i_addr_rom[  269] = 'h000002a8; 	    d_addr_rom[  269] = 'h00000a88; 	    wdata_rom[  269] = 'h255f47bb; 	    wvalid_rom[  269] = 0; 
    i_addr_rom[  270] = 'h0000051c; 	    d_addr_rom[  270] = 'h0000093c; 	    wdata_rom[  270] = 'h1118149e; 	    wvalid_rom[  270] = 1; 
    i_addr_rom[  271] = 'h000000ec; 	    d_addr_rom[  271] = 'h00000e94; 	    wdata_rom[  271] = 'h04aafe83; 	    wvalid_rom[  271] = 1; 
    i_addr_rom[  272] = 'h0000054c; 	    d_addr_rom[  272] = 'h00000c44; 	    wdata_rom[  272] = 'hd49eaf5a; 	    wvalid_rom[  272] = 0; 
    i_addr_rom[  273] = 'h00000184; 	    d_addr_rom[  273] = 'h00000c20; 	    wdata_rom[  273] = 'h41229175; 	    wvalid_rom[  273] = 0; 
    i_addr_rom[  274] = 'h00000628; 	    d_addr_rom[  274] = 'h00000938; 	    wdata_rom[  274] = 'h9edc3bfd; 	    wvalid_rom[  274] = 1; 
    i_addr_rom[  275] = 'h0000051c; 	    d_addr_rom[  275] = 'h00000900; 	    wdata_rom[  275] = 'h2ca391c2; 	    wvalid_rom[  275] = 0; 
    i_addr_rom[  276] = 'h000006b8; 	    d_addr_rom[  276] = 'h00000ef0; 	    wdata_rom[  276] = 'h16c675e1; 	    wvalid_rom[  276] = 1; 
    i_addr_rom[  277] = 'h000007c8; 	    d_addr_rom[  277] = 'h00000a64; 	    wdata_rom[  277] = 'h43fafb53; 	    wvalid_rom[  277] = 0; 
    i_addr_rom[  278] = 'h0000022c; 	    d_addr_rom[  278] = 'h00000a6c; 	    wdata_rom[  278] = 'heb11844e; 	    wvalid_rom[  278] = 1; 
    i_addr_rom[  279] = 'h00000424; 	    d_addr_rom[  279] = 'h00000d70; 	    wdata_rom[  279] = 'hccd3fbe7; 	    wvalid_rom[  279] = 1; 
    i_addr_rom[  280] = 'h000001b0; 	    d_addr_rom[  280] = 'h00000ba8; 	    wdata_rom[  280] = 'h132b41f2; 	    wvalid_rom[  280] = 0; 
    i_addr_rom[  281] = 'h000001f4; 	    d_addr_rom[  281] = 'h00000f20; 	    wdata_rom[  281] = 'h74fa5fb8; 	    wvalid_rom[  281] = 1; 
    i_addr_rom[  282] = 'h000007cc; 	    d_addr_rom[  282] = 'h00000d0c; 	    wdata_rom[  282] = 'h83feb940; 	    wvalid_rom[  282] = 0; 
    i_addr_rom[  283] = 'h0000074c; 	    d_addr_rom[  283] = 'h00000cd4; 	    wdata_rom[  283] = 'h87b6e9df; 	    wvalid_rom[  283] = 1; 
    i_addr_rom[  284] = 'h00000598; 	    d_addr_rom[  284] = 'h0000085c; 	    wdata_rom[  284] = 'h8bcd94bb; 	    wvalid_rom[  284] = 1; 
    i_addr_rom[  285] = 'h00000508; 	    d_addr_rom[  285] = 'h00000d7c; 	    wdata_rom[  285] = 'hb5f45719; 	    wvalid_rom[  285] = 0; 
    i_addr_rom[  286] = 'h000004bc; 	    d_addr_rom[  286] = 'h00000f08; 	    wdata_rom[  286] = 'h6b74954d; 	    wvalid_rom[  286] = 1; 
    i_addr_rom[  287] = 'h0000019c; 	    d_addr_rom[  287] = 'h00000d88; 	    wdata_rom[  287] = 'h5d3ff1f8; 	    wvalid_rom[  287] = 1; 
    i_addr_rom[  288] = 'h000002b4; 	    d_addr_rom[  288] = 'h000009ac; 	    wdata_rom[  288] = 'h0d890f51; 	    wvalid_rom[  288] = 1; 
    i_addr_rom[  289] = 'h0000065c; 	    d_addr_rom[  289] = 'h00000cd8; 	    wdata_rom[  289] = 'he013fb46; 	    wvalid_rom[  289] = 0; 
    i_addr_rom[  290] = 'h0000018c; 	    d_addr_rom[  290] = 'h00000af8; 	    wdata_rom[  290] = 'h3222e1dd; 	    wvalid_rom[  290] = 1; 
    i_addr_rom[  291] = 'h00000350; 	    d_addr_rom[  291] = 'h00000b5c; 	    wdata_rom[  291] = 'h756564b5; 	    wvalid_rom[  291] = 0; 
    i_addr_rom[  292] = 'h000001a8; 	    d_addr_rom[  292] = 'h00000920; 	    wdata_rom[  292] = 'h892d5ee9; 	    wvalid_rom[  292] = 1; 
    i_addr_rom[  293] = 'h00000524; 	    d_addr_rom[  293] = 'h0000099c; 	    wdata_rom[  293] = 'hb7c162b8; 	    wvalid_rom[  293] = 1; 
    i_addr_rom[  294] = 'h00000350; 	    d_addr_rom[  294] = 'h00000f94; 	    wdata_rom[  294] = 'h950c48b9; 	    wvalid_rom[  294] = 1; 
    i_addr_rom[  295] = 'h000000b4; 	    d_addr_rom[  295] = 'h00000ad0; 	    wdata_rom[  295] = 'h6d5ea936; 	    wvalid_rom[  295] = 1; 
    i_addr_rom[  296] = 'h000001f8; 	    d_addr_rom[  296] = 'h00000ad8; 	    wdata_rom[  296] = 'h220ff094; 	    wvalid_rom[  296] = 0; 
    i_addr_rom[  297] = 'h000004c8; 	    d_addr_rom[  297] = 'h00000ee8; 	    wdata_rom[  297] = 'h024ef9cc; 	    wvalid_rom[  297] = 0; 
    i_addr_rom[  298] = 'h00000458; 	    d_addr_rom[  298] = 'h00000a5c; 	    wdata_rom[  298] = 'h77e0e453; 	    wvalid_rom[  298] = 1; 
    i_addr_rom[  299] = 'h000006d4; 	    d_addr_rom[  299] = 'h00000acc; 	    wdata_rom[  299] = 'hda63c358; 	    wvalid_rom[  299] = 1; 
    i_addr_rom[  300] = 'h00000680; 	    d_addr_rom[  300] = 'h00000d2c; 	    wdata_rom[  300] = 'h528e01d5; 	    wvalid_rom[  300] = 1; 
    i_addr_rom[  301] = 'h000004fc; 	    d_addr_rom[  301] = 'h00000fd0; 	    wdata_rom[  301] = 'h38cc812d; 	    wvalid_rom[  301] = 0; 
    i_addr_rom[  302] = 'h00000574; 	    d_addr_rom[  302] = 'h00000918; 	    wdata_rom[  302] = 'hcd356549; 	    wvalid_rom[  302] = 1; 
    i_addr_rom[  303] = 'h0000018c; 	    d_addr_rom[  303] = 'h00000954; 	    wdata_rom[  303] = 'h7fad8564; 	    wvalid_rom[  303] = 0; 
    i_addr_rom[  304] = 'h0000062c; 	    d_addr_rom[  304] = 'h00000c64; 	    wdata_rom[  304] = 'ha70a25b3; 	    wvalid_rom[  304] = 0; 
    i_addr_rom[  305] = 'h000006b8; 	    d_addr_rom[  305] = 'h00000a40; 	    wdata_rom[  305] = 'ha7de6433; 	    wvalid_rom[  305] = 0; 
    i_addr_rom[  306] = 'h000003d4; 	    d_addr_rom[  306] = 'h00000ae8; 	    wdata_rom[  306] = 'h4d0bad27; 	    wvalid_rom[  306] = 0; 
    i_addr_rom[  307] = 'h00000470; 	    d_addr_rom[  307] = 'h00000888; 	    wdata_rom[  307] = 'h6cd5d160; 	    wvalid_rom[  307] = 0; 
    i_addr_rom[  308] = 'h00000104; 	    d_addr_rom[  308] = 'h00000fb4; 	    wdata_rom[  308] = 'h473b1627; 	    wvalid_rom[  308] = 1; 
    i_addr_rom[  309] = 'h0000032c; 	    d_addr_rom[  309] = 'h00000f40; 	    wdata_rom[  309] = 'h0148fabe; 	    wvalid_rom[  309] = 0; 
    i_addr_rom[  310] = 'h000000c4; 	    d_addr_rom[  310] = 'h00000818; 	    wdata_rom[  310] = 'h6fd4c7a5; 	    wvalid_rom[  310] = 0; 
    i_addr_rom[  311] = 'h000001c8; 	    d_addr_rom[  311] = 'h00000ba0; 	    wdata_rom[  311] = 'hbaa3ee5b; 	    wvalid_rom[  311] = 1; 
    i_addr_rom[  312] = 'h0000068c; 	    d_addr_rom[  312] = 'h00000c58; 	    wdata_rom[  312] = 'h6c94ade4; 	    wvalid_rom[  312] = 0; 
    i_addr_rom[  313] = 'h00000474; 	    d_addr_rom[  313] = 'h00000ea0; 	    wdata_rom[  313] = 'h7d7c4adf; 	    wvalid_rom[  313] = 0; 
    i_addr_rom[  314] = 'h000005e0; 	    d_addr_rom[  314] = 'h00000acc; 	    wdata_rom[  314] = 'h48bb7637; 	    wvalid_rom[  314] = 1; 
    i_addr_rom[  315] = 'h00000498; 	    d_addr_rom[  315] = 'h00000d1c; 	    wdata_rom[  315] = 'h4bbbe52d; 	    wvalid_rom[  315] = 0; 
    i_addr_rom[  316] = 'h00000768; 	    d_addr_rom[  316] = 'h00000c28; 	    wdata_rom[  316] = 'ha6209f49; 	    wvalid_rom[  316] = 1; 
    i_addr_rom[  317] = 'h000007cc; 	    d_addr_rom[  317] = 'h00000c68; 	    wdata_rom[  317] = 'hbaed18c8; 	    wvalid_rom[  317] = 0; 
    i_addr_rom[  318] = 'h00000414; 	    d_addr_rom[  318] = 'h00000c0c; 	    wdata_rom[  318] = 'hd737b749; 	    wvalid_rom[  318] = 1; 
    i_addr_rom[  319] = 'h00000600; 	    d_addr_rom[  319] = 'h00000cf0; 	    wdata_rom[  319] = 'ha63fc8cc; 	    wvalid_rom[  319] = 1; 
    i_addr_rom[  320] = 'h000001cc; 	    d_addr_rom[  320] = 'h00000c34; 	    wdata_rom[  320] = 'h029943f0; 	    wvalid_rom[  320] = 1; 
    i_addr_rom[  321] = 'h0000041c; 	    d_addr_rom[  321] = 'h00000f4c; 	    wdata_rom[  321] = 'hc04afb32; 	    wvalid_rom[  321] = 1; 
    i_addr_rom[  322] = 'h000004b0; 	    d_addr_rom[  322] = 'h00000ff0; 	    wdata_rom[  322] = 'h18a07f8a; 	    wvalid_rom[  322] = 1; 
    i_addr_rom[  323] = 'h0000031c; 	    d_addr_rom[  323] = 'h00000ecc; 	    wdata_rom[  323] = 'he6d2d82d; 	    wvalid_rom[  323] = 0; 
    i_addr_rom[  324] = 'h000007d4; 	    d_addr_rom[  324] = 'h00000830; 	    wdata_rom[  324] = 'h691a43e5; 	    wvalid_rom[  324] = 0; 
    i_addr_rom[  325] = 'h000006bc; 	    d_addr_rom[  325] = 'h000009b8; 	    wdata_rom[  325] = 'hc3fed1e5; 	    wvalid_rom[  325] = 1; 
    i_addr_rom[  326] = 'h000003e4; 	    d_addr_rom[  326] = 'h00000954; 	    wdata_rom[  326] = 'hf3008ca8; 	    wvalid_rom[  326] = 1; 
    i_addr_rom[  327] = 'h000003a0; 	    d_addr_rom[  327] = 'h00000fc4; 	    wdata_rom[  327] = 'h2bbf7741; 	    wvalid_rom[  327] = 1; 
    i_addr_rom[  328] = 'h00000584; 	    d_addr_rom[  328] = 'h00000ad0; 	    wdata_rom[  328] = 'hdbcb296f; 	    wvalid_rom[  328] = 1; 
    i_addr_rom[  329] = 'h000000fc; 	    d_addr_rom[  329] = 'h00000bdc; 	    wdata_rom[  329] = 'h7322f856; 	    wvalid_rom[  329] = 1; 
    i_addr_rom[  330] = 'h000003b8; 	    d_addr_rom[  330] = 'h0000098c; 	    wdata_rom[  330] = 'h955a5a77; 	    wvalid_rom[  330] = 1; 
    i_addr_rom[  331] = 'h00000384; 	    d_addr_rom[  331] = 'h00000810; 	    wdata_rom[  331] = 'h2c33bcd9; 	    wvalid_rom[  331] = 0; 
    i_addr_rom[  332] = 'h00000284; 	    d_addr_rom[  332] = 'h00000800; 	    wdata_rom[  332] = 'hde0c08be; 	    wvalid_rom[  332] = 0; 
    i_addr_rom[  333] = 'h000002d0; 	    d_addr_rom[  333] = 'h00000d9c; 	    wdata_rom[  333] = 'hcb286eaa; 	    wvalid_rom[  333] = 0; 
    i_addr_rom[  334] = 'h000006e4; 	    d_addr_rom[  334] = 'h00000d30; 	    wdata_rom[  334] = 'hdc0a2c66; 	    wvalid_rom[  334] = 0; 
    i_addr_rom[  335] = 'h0000049c; 	    d_addr_rom[  335] = 'h00000b20; 	    wdata_rom[  335] = 'h6d2ec712; 	    wvalid_rom[  335] = 0; 
    i_addr_rom[  336] = 'h000005e0; 	    d_addr_rom[  336] = 'h00000d64; 	    wdata_rom[  336] = 'h0f6fe760; 	    wvalid_rom[  336] = 0; 
    i_addr_rom[  337] = 'h00000144; 	    d_addr_rom[  337] = 'h000008bc; 	    wdata_rom[  337] = 'h62d87ed6; 	    wvalid_rom[  337] = 1; 
    i_addr_rom[  338] = 'h0000047c; 	    d_addr_rom[  338] = 'h00000b1c; 	    wdata_rom[  338] = 'h68f5d9fa; 	    wvalid_rom[  338] = 0; 
    i_addr_rom[  339] = 'h00000378; 	    d_addr_rom[  339] = 'h00000d48; 	    wdata_rom[  339] = 'h33b375ab; 	    wvalid_rom[  339] = 1; 
    i_addr_rom[  340] = 'h000004f0; 	    d_addr_rom[  340] = 'h000009b8; 	    wdata_rom[  340] = 'h24376575; 	    wvalid_rom[  340] = 0; 
    i_addr_rom[  341] = 'h00000274; 	    d_addr_rom[  341] = 'h00000f94; 	    wdata_rom[  341] = 'h2102ea9a; 	    wvalid_rom[  341] = 0; 
    i_addr_rom[  342] = 'h000004ec; 	    d_addr_rom[  342] = 'h00000aa0; 	    wdata_rom[  342] = 'h4a730b04; 	    wvalid_rom[  342] = 0; 
    i_addr_rom[  343] = 'h000002b8; 	    d_addr_rom[  343] = 'h00000bbc; 	    wdata_rom[  343] = 'h69315ba0; 	    wvalid_rom[  343] = 1; 
    i_addr_rom[  344] = 'h000002a0; 	    d_addr_rom[  344] = 'h00000af4; 	    wdata_rom[  344] = 'h9b76fae9; 	    wvalid_rom[  344] = 1; 
    i_addr_rom[  345] = 'h00000730; 	    d_addr_rom[  345] = 'h00000cfc; 	    wdata_rom[  345] = 'h675690ca; 	    wvalid_rom[  345] = 0; 
    i_addr_rom[  346] = 'h00000794; 	    d_addr_rom[  346] = 'h00000e40; 	    wdata_rom[  346] = 'h91a8ff5d; 	    wvalid_rom[  346] = 0; 
    i_addr_rom[  347] = 'h000004e8; 	    d_addr_rom[  347] = 'h000009b0; 	    wdata_rom[  347] = 'hc3417fce; 	    wvalid_rom[  347] = 1; 
    i_addr_rom[  348] = 'h00000418; 	    d_addr_rom[  348] = 'h00000e50; 	    wdata_rom[  348] = 'hffbc00e7; 	    wvalid_rom[  348] = 0; 
    i_addr_rom[  349] = 'h000001f0; 	    d_addr_rom[  349] = 'h000009d8; 	    wdata_rom[  349] = 'h1d656b0a; 	    wvalid_rom[  349] = 0; 
    i_addr_rom[  350] = 'h000006a0; 	    d_addr_rom[  350] = 'h00000ba8; 	    wdata_rom[  350] = 'h4526e956; 	    wvalid_rom[  350] = 0; 
    i_addr_rom[  351] = 'h00000130; 	    d_addr_rom[  351] = 'h00000eac; 	    wdata_rom[  351] = 'h56b71c4c; 	    wvalid_rom[  351] = 1; 
    i_addr_rom[  352] = 'h00000618; 	    d_addr_rom[  352] = 'h00000c74; 	    wdata_rom[  352] = 'h54967ffe; 	    wvalid_rom[  352] = 1; 
    i_addr_rom[  353] = 'h000001f8; 	    d_addr_rom[  353] = 'h00000aac; 	    wdata_rom[  353] = 'h11e0a9e1; 	    wvalid_rom[  353] = 0; 
    i_addr_rom[  354] = 'h00000768; 	    d_addr_rom[  354] = 'h00000e54; 	    wdata_rom[  354] = 'h73ee62ea; 	    wvalid_rom[  354] = 1; 
    i_addr_rom[  355] = 'h00000060; 	    d_addr_rom[  355] = 'h000009cc; 	    wdata_rom[  355] = 'h362a2164; 	    wvalid_rom[  355] = 0; 
    i_addr_rom[  356] = 'h00000160; 	    d_addr_rom[  356] = 'h00000b0c; 	    wdata_rom[  356] = 'hd3fd4f0c; 	    wvalid_rom[  356] = 0; 
    i_addr_rom[  357] = 'h00000570; 	    d_addr_rom[  357] = 'h00000c9c; 	    wdata_rom[  357] = 'h420163e3; 	    wvalid_rom[  357] = 1; 
    i_addr_rom[  358] = 'h000006f0; 	    d_addr_rom[  358] = 'h00000920; 	    wdata_rom[  358] = 'h74004e3d; 	    wvalid_rom[  358] = 0; 
    i_addr_rom[  359] = 'h000007f8; 	    d_addr_rom[  359] = 'h0000093c; 	    wdata_rom[  359] = 'hcdf420e5; 	    wvalid_rom[  359] = 1; 
    i_addr_rom[  360] = 'h00000148; 	    d_addr_rom[  360] = 'h00000a34; 	    wdata_rom[  360] = 'he11e5aaf; 	    wvalid_rom[  360] = 1; 
    i_addr_rom[  361] = 'h000007e8; 	    d_addr_rom[  361] = 'h00000ccc; 	    wdata_rom[  361] = 'h81f0f809; 	    wvalid_rom[  361] = 1; 
    i_addr_rom[  362] = 'h00000138; 	    d_addr_rom[  362] = 'h00000efc; 	    wdata_rom[  362] = 'h7ab2e575; 	    wvalid_rom[  362] = 0; 
    i_addr_rom[  363] = 'h00000484; 	    d_addr_rom[  363] = 'h00000c20; 	    wdata_rom[  363] = 'h67bd215a; 	    wvalid_rom[  363] = 1; 
    i_addr_rom[  364] = 'h000003f8; 	    d_addr_rom[  364] = 'h00000be8; 	    wdata_rom[  364] = 'h8aa5a071; 	    wvalid_rom[  364] = 1; 
    i_addr_rom[  365] = 'h00000378; 	    d_addr_rom[  365] = 'h00000d6c; 	    wdata_rom[  365] = 'h8042d8de; 	    wvalid_rom[  365] = 1; 
    i_addr_rom[  366] = 'h00000604; 	    d_addr_rom[  366] = 'h00000b9c; 	    wdata_rom[  366] = 'h3c83b178; 	    wvalid_rom[  366] = 0; 
    i_addr_rom[  367] = 'h00000650; 	    d_addr_rom[  367] = 'h00000a2c; 	    wdata_rom[  367] = 'h22006692; 	    wvalid_rom[  367] = 1; 
    i_addr_rom[  368] = 'h000004a0; 	    d_addr_rom[  368] = 'h00000b60; 	    wdata_rom[  368] = 'h806e7228; 	    wvalid_rom[  368] = 0; 
    i_addr_rom[  369] = 'h0000025c; 	    d_addr_rom[  369] = 'h00000dc4; 	    wdata_rom[  369] = 'hb2ec1674; 	    wvalid_rom[  369] = 0; 
    i_addr_rom[  370] = 'h00000628; 	    d_addr_rom[  370] = 'h00000a9c; 	    wdata_rom[  370] = 'h854a4dc8; 	    wvalid_rom[  370] = 0; 
    i_addr_rom[  371] = 'h00000370; 	    d_addr_rom[  371] = 'h0000094c; 	    wdata_rom[  371] = 'hf108e903; 	    wvalid_rom[  371] = 0; 
    i_addr_rom[  372] = 'h0000018c; 	    d_addr_rom[  372] = 'h00000eec; 	    wdata_rom[  372] = 'h5c7435a5; 	    wvalid_rom[  372] = 1; 
    i_addr_rom[  373] = 'h0000047c; 	    d_addr_rom[  373] = 'h00000984; 	    wdata_rom[  373] = 'ha2626e95; 	    wvalid_rom[  373] = 1; 
    i_addr_rom[  374] = 'h000005c0; 	    d_addr_rom[  374] = 'h00000ff4; 	    wdata_rom[  374] = 'h6c52c30f; 	    wvalid_rom[  374] = 1; 
    i_addr_rom[  375] = 'h000003e0; 	    d_addr_rom[  375] = 'h00000ef8; 	    wdata_rom[  375] = 'h59b06d58; 	    wvalid_rom[  375] = 0; 
    i_addr_rom[  376] = 'h000006c8; 	    d_addr_rom[  376] = 'h00000f70; 	    wdata_rom[  376] = 'h96c27098; 	    wvalid_rom[  376] = 0; 
    i_addr_rom[  377] = 'h00000118; 	    d_addr_rom[  377] = 'h000008d4; 	    wdata_rom[  377] = 'hc6b8d9d4; 	    wvalid_rom[  377] = 1; 
    i_addr_rom[  378] = 'h00000688; 	    d_addr_rom[  378] = 'h00000a34; 	    wdata_rom[  378] = 'h72839828; 	    wvalid_rom[  378] = 0; 
    i_addr_rom[  379] = 'h00000290; 	    d_addr_rom[  379] = 'h00000f2c; 	    wdata_rom[  379] = 'h3cd2ada9; 	    wvalid_rom[  379] = 0; 
    i_addr_rom[  380] = 'h00000720; 	    d_addr_rom[  380] = 'h00000a4c; 	    wdata_rom[  380] = 'h37ff4dcf; 	    wvalid_rom[  380] = 0; 
    i_addr_rom[  381] = 'h000002d0; 	    d_addr_rom[  381] = 'h000009a4; 	    wdata_rom[  381] = 'he0c08215; 	    wvalid_rom[  381] = 0; 
    i_addr_rom[  382] = 'h0000009c; 	    d_addr_rom[  382] = 'h00000b54; 	    wdata_rom[  382] = 'h63188d8e; 	    wvalid_rom[  382] = 0; 
    i_addr_rom[  383] = 'h00000334; 	    d_addr_rom[  383] = 'h00000a64; 	    wdata_rom[  383] = 'h0b85e8b2; 	    wvalid_rom[  383] = 0; 
    i_addr_rom[  384] = 'h0000062c; 	    d_addr_rom[  384] = 'h00000b24; 	    wdata_rom[  384] = 'h6ea0447e; 	    wvalid_rom[  384] = 0; 
    i_addr_rom[  385] = 'h00000678; 	    d_addr_rom[  385] = 'h00000924; 	    wdata_rom[  385] = 'hf8890620; 	    wvalid_rom[  385] = 0; 
    i_addr_rom[  386] = 'h0000059c; 	    d_addr_rom[  386] = 'h00000f6c; 	    wdata_rom[  386] = 'h9e3d2928; 	    wvalid_rom[  386] = 0; 
    i_addr_rom[  387] = 'h000007c4; 	    d_addr_rom[  387] = 'h00000ab8; 	    wdata_rom[  387] = 'he9cfafee; 	    wvalid_rom[  387] = 0; 
    i_addr_rom[  388] = 'h00000584; 	    d_addr_rom[  388] = 'h00000fc4; 	    wdata_rom[  388] = 'h63b6f382; 	    wvalid_rom[  388] = 1; 
    i_addr_rom[  389] = 'h0000041c; 	    d_addr_rom[  389] = 'h00000ffc; 	    wdata_rom[  389] = 'h0a892165; 	    wvalid_rom[  389] = 0; 
    i_addr_rom[  390] = 'h00000308; 	    d_addr_rom[  390] = 'h00000c20; 	    wdata_rom[  390] = 'h7353bc3f; 	    wvalid_rom[  390] = 1; 
    i_addr_rom[  391] = 'h000003bc; 	    d_addr_rom[  391] = 'h00000e34; 	    wdata_rom[  391] = 'h58d4ccfd; 	    wvalid_rom[  391] = 1; 
    i_addr_rom[  392] = 'h00000468; 	    d_addr_rom[  392] = 'h00000fe0; 	    wdata_rom[  392] = 'hdb48f66d; 	    wvalid_rom[  392] = 0; 
    i_addr_rom[  393] = 'h00000460; 	    d_addr_rom[  393] = 'h00000838; 	    wdata_rom[  393] = 'hab90e523; 	    wvalid_rom[  393] = 1; 
    i_addr_rom[  394] = 'h000000ec; 	    d_addr_rom[  394] = 'h00000ea4; 	    wdata_rom[  394] = 'h0bdae1f5; 	    wvalid_rom[  394] = 0; 
    i_addr_rom[  395] = 'h00000434; 	    d_addr_rom[  395] = 'h00000820; 	    wdata_rom[  395] = 'h98845da1; 	    wvalid_rom[  395] = 0; 
    i_addr_rom[  396] = 'h000002d8; 	    d_addr_rom[  396] = 'h00000c80; 	    wdata_rom[  396] = 'h52074d31; 	    wvalid_rom[  396] = 1; 
    i_addr_rom[  397] = 'h0000072c; 	    d_addr_rom[  397] = 'h00000d3c; 	    wdata_rom[  397] = 'h5cfe2e3e; 	    wvalid_rom[  397] = 1; 
    i_addr_rom[  398] = 'h000000cc; 	    d_addr_rom[  398] = 'h00000c44; 	    wdata_rom[  398] = 'hf4a55c13; 	    wvalid_rom[  398] = 1; 
    i_addr_rom[  399] = 'h00000120; 	    d_addr_rom[  399] = 'h00000de4; 	    wdata_rom[  399] = 'h35cf1edb; 	    wvalid_rom[  399] = 0; 
    i_addr_rom[  400] = 'h000005f0; 	    d_addr_rom[  400] = 'h00000a90; 	    wdata_rom[  400] = 'h9552b863; 	    wvalid_rom[  400] = 0; 
    i_addr_rom[  401] = 'h00000794; 	    d_addr_rom[  401] = 'h000009f0; 	    wdata_rom[  401] = 'h216607d6; 	    wvalid_rom[  401] = 0; 
    i_addr_rom[  402] = 'h00000258; 	    d_addr_rom[  402] = 'h00000ee8; 	    wdata_rom[  402] = 'hef2c5626; 	    wvalid_rom[  402] = 1; 
    i_addr_rom[  403] = 'h000000a0; 	    d_addr_rom[  403] = 'h00000d08; 	    wdata_rom[  403] = 'h4010864c; 	    wvalid_rom[  403] = 1; 
    i_addr_rom[  404] = 'h000002d8; 	    d_addr_rom[  404] = 'h000009e4; 	    wdata_rom[  404] = 'hd90f07c1; 	    wvalid_rom[  404] = 0; 
    i_addr_rom[  405] = 'h00000670; 	    d_addr_rom[  405] = 'h00000efc; 	    wdata_rom[  405] = 'ha7d9c3d9; 	    wvalid_rom[  405] = 0; 
    i_addr_rom[  406] = 'h000007e4; 	    d_addr_rom[  406] = 'h00000928; 	    wdata_rom[  406] = 'h7fd8d5e5; 	    wvalid_rom[  406] = 1; 
    i_addr_rom[  407] = 'h000002f4; 	    d_addr_rom[  407] = 'h00000f08; 	    wdata_rom[  407] = 'h5fd63b74; 	    wvalid_rom[  407] = 1; 
    i_addr_rom[  408] = 'h00000034; 	    d_addr_rom[  408] = 'h000009e4; 	    wdata_rom[  408] = 'h2549db0f; 	    wvalid_rom[  408] = 1; 
    i_addr_rom[  409] = 'h00000208; 	    d_addr_rom[  409] = 'h00000fc0; 	    wdata_rom[  409] = 'h4e517647; 	    wvalid_rom[  409] = 0; 
    i_addr_rom[  410] = 'h00000738; 	    d_addr_rom[  410] = 'h00000c14; 	    wdata_rom[  410] = 'hfac416da; 	    wvalid_rom[  410] = 1; 
    i_addr_rom[  411] = 'h00000504; 	    d_addr_rom[  411] = 'h00000d4c; 	    wdata_rom[  411] = 'h50a03b75; 	    wvalid_rom[  411] = 1; 
    i_addr_rom[  412] = 'h000004c4; 	    d_addr_rom[  412] = 'h00000e10; 	    wdata_rom[  412] = 'h2b775e7e; 	    wvalid_rom[  412] = 0; 
    i_addr_rom[  413] = 'h000007a8; 	    d_addr_rom[  413] = 'h00000e58; 	    wdata_rom[  413] = 'hc9de9ec9; 	    wvalid_rom[  413] = 1; 
    i_addr_rom[  414] = 'h000007d4; 	    d_addr_rom[  414] = 'h00000ac0; 	    wdata_rom[  414] = 'hd0c145de; 	    wvalid_rom[  414] = 1; 
    i_addr_rom[  415] = 'h00000360; 	    d_addr_rom[  415] = 'h000008e8; 	    wdata_rom[  415] = 'hed9787e7; 	    wvalid_rom[  415] = 1; 
    i_addr_rom[  416] = 'h00000460; 	    d_addr_rom[  416] = 'h00000b64; 	    wdata_rom[  416] = 'habb17763; 	    wvalid_rom[  416] = 0; 
    i_addr_rom[  417] = 'h00000090; 	    d_addr_rom[  417] = 'h000009d8; 	    wdata_rom[  417] = 'h756b32ba; 	    wvalid_rom[  417] = 1; 
    i_addr_rom[  418] = 'h0000079c; 	    d_addr_rom[  418] = 'h00000c40; 	    wdata_rom[  418] = 'h17dad1ed; 	    wvalid_rom[  418] = 0; 
    i_addr_rom[  419] = 'h000007fc; 	    d_addr_rom[  419] = 'h00000cb0; 	    wdata_rom[  419] = 'haa624248; 	    wvalid_rom[  419] = 1; 
    i_addr_rom[  420] = 'h00000330; 	    d_addr_rom[  420] = 'h00000cd4; 	    wdata_rom[  420] = 'hc5cb33b4; 	    wvalid_rom[  420] = 1; 
    i_addr_rom[  421] = 'h00000470; 	    d_addr_rom[  421] = 'h00000904; 	    wdata_rom[  421] = 'hbe4b624f; 	    wvalid_rom[  421] = 0; 
    i_addr_rom[  422] = 'h00000128; 	    d_addr_rom[  422] = 'h00000fe4; 	    wdata_rom[  422] = 'h2e8c1efc; 	    wvalid_rom[  422] = 1; 
    i_addr_rom[  423] = 'h000007c0; 	    d_addr_rom[  423] = 'h00000ff4; 	    wdata_rom[  423] = 'h617db5ed; 	    wvalid_rom[  423] = 1; 
    i_addr_rom[  424] = 'h000001f4; 	    d_addr_rom[  424] = 'h00000d74; 	    wdata_rom[  424] = 'h316310ba; 	    wvalid_rom[  424] = 1; 
    i_addr_rom[  425] = 'h00000638; 	    d_addr_rom[  425] = 'h00000c58; 	    wdata_rom[  425] = 'h3b726e30; 	    wvalid_rom[  425] = 1; 
    i_addr_rom[  426] = 'h0000070c; 	    d_addr_rom[  426] = 'h00000e20; 	    wdata_rom[  426] = 'h31af39b9; 	    wvalid_rom[  426] = 1; 
    i_addr_rom[  427] = 'h00000554; 	    d_addr_rom[  427] = 'h00000994; 	    wdata_rom[  427] = 'he34bd20d; 	    wvalid_rom[  427] = 1; 
    i_addr_rom[  428] = 'h000000fc; 	    d_addr_rom[  428] = 'h00000ccc; 	    wdata_rom[  428] = 'h2e99f1f7; 	    wvalid_rom[  428] = 1; 
    i_addr_rom[  429] = 'h0000053c; 	    d_addr_rom[  429] = 'h00000a74; 	    wdata_rom[  429] = 'h1fef3fcf; 	    wvalid_rom[  429] = 0; 
    i_addr_rom[  430] = 'h000003e8; 	    d_addr_rom[  430] = 'h00000b68; 	    wdata_rom[  430] = 'h3e89c667; 	    wvalid_rom[  430] = 1; 
    i_addr_rom[  431] = 'h00000774; 	    d_addr_rom[  431] = 'h00000de4; 	    wdata_rom[  431] = 'hee0caa8f; 	    wvalid_rom[  431] = 0; 
    i_addr_rom[  432] = 'h00000368; 	    d_addr_rom[  432] = 'h00000fdc; 	    wdata_rom[  432] = 'h25cac425; 	    wvalid_rom[  432] = 1; 
    i_addr_rom[  433] = 'h00000520; 	    d_addr_rom[  433] = 'h00000864; 	    wdata_rom[  433] = 'h97a28278; 	    wvalid_rom[  433] = 1; 
    i_addr_rom[  434] = 'h000003e8; 	    d_addr_rom[  434] = 'h00000c3c; 	    wdata_rom[  434] = 'h7137457b; 	    wvalid_rom[  434] = 0; 
    i_addr_rom[  435] = 'h000002bc; 	    d_addr_rom[  435] = 'h00000e00; 	    wdata_rom[  435] = 'ha0967c66; 	    wvalid_rom[  435] = 0; 
    i_addr_rom[  436] = 'h0000057c; 	    d_addr_rom[  436] = 'h000008e4; 	    wdata_rom[  436] = 'he33540f6; 	    wvalid_rom[  436] = 0; 
    i_addr_rom[  437] = 'h000002e0; 	    d_addr_rom[  437] = 'h000009f0; 	    wdata_rom[  437] = 'h976edf44; 	    wvalid_rom[  437] = 0; 
    i_addr_rom[  438] = 'h0000037c; 	    d_addr_rom[  438] = 'h00000844; 	    wdata_rom[  438] = 'hdc066570; 	    wvalid_rom[  438] = 1; 
    i_addr_rom[  439] = 'h00000534; 	    d_addr_rom[  439] = 'h00000ba4; 	    wdata_rom[  439] = 'h9d239c86; 	    wvalid_rom[  439] = 1; 
    i_addr_rom[  440] = 'h00000198; 	    d_addr_rom[  440] = 'h00000a60; 	    wdata_rom[  440] = 'h8eaf3cb1; 	    wvalid_rom[  440] = 1; 
    i_addr_rom[  441] = 'h00000748; 	    d_addr_rom[  441] = 'h00000ae8; 	    wdata_rom[  441] = 'hce3356ce; 	    wvalid_rom[  441] = 0; 
    i_addr_rom[  442] = 'h00000618; 	    d_addr_rom[  442] = 'h00000c20; 	    wdata_rom[  442] = 'h57603941; 	    wvalid_rom[  442] = 1; 
    i_addr_rom[  443] = 'h00000000; 	    d_addr_rom[  443] = 'h00000d08; 	    wdata_rom[  443] = 'he0cba9e4; 	    wvalid_rom[  443] = 0; 
    i_addr_rom[  444] = 'h00000390; 	    d_addr_rom[  444] = 'h0000098c; 	    wdata_rom[  444] = 'h07004c70; 	    wvalid_rom[  444] = 0; 
    i_addr_rom[  445] = 'h00000138; 	    d_addr_rom[  445] = 'h00000abc; 	    wdata_rom[  445] = 'hbb0be6da; 	    wvalid_rom[  445] = 1; 
    i_addr_rom[  446] = 'h00000694; 	    d_addr_rom[  446] = 'h00000d54; 	    wdata_rom[  446] = 'ha75d5934; 	    wvalid_rom[  446] = 1; 
    i_addr_rom[  447] = 'h000001bc; 	    d_addr_rom[  447] = 'h00000a10; 	    wdata_rom[  447] = 'hf9a9bd5b; 	    wvalid_rom[  447] = 0; 
    i_addr_rom[  448] = 'h000007bc; 	    d_addr_rom[  448] = 'h00000f64; 	    wdata_rom[  448] = 'hba55eceb; 	    wvalid_rom[  448] = 0; 
    i_addr_rom[  449] = 'h0000019c; 	    d_addr_rom[  449] = 'h00000ce0; 	    wdata_rom[  449] = 'hb22b4b07; 	    wvalid_rom[  449] = 1; 
    i_addr_rom[  450] = 'h0000046c; 	    d_addr_rom[  450] = 'h00000ff8; 	    wdata_rom[  450] = 'h7b60c85e; 	    wvalid_rom[  450] = 1; 
    i_addr_rom[  451] = 'h00000574; 	    d_addr_rom[  451] = 'h0000099c; 	    wdata_rom[  451] = 'hf24b1dfa; 	    wvalid_rom[  451] = 1; 
    i_addr_rom[  452] = 'h00000650; 	    d_addr_rom[  452] = 'h0000087c; 	    wdata_rom[  452] = 'h4caceb77; 	    wvalid_rom[  452] = 1; 
    i_addr_rom[  453] = 'h000003c0; 	    d_addr_rom[  453] = 'h00000840; 	    wdata_rom[  453] = 'h13eadf3b; 	    wvalid_rom[  453] = 0; 
    i_addr_rom[  454] = 'h0000055c; 	    d_addr_rom[  454] = 'h00000ed4; 	    wdata_rom[  454] = 'heb3b228e; 	    wvalid_rom[  454] = 0; 
    i_addr_rom[  455] = 'h00000170; 	    d_addr_rom[  455] = 'h00000844; 	    wdata_rom[  455] = 'h1a2930e9; 	    wvalid_rom[  455] = 0; 
    i_addr_rom[  456] = 'h00000068; 	    d_addr_rom[  456] = 'h00000bb8; 	    wdata_rom[  456] = 'h85d22a41; 	    wvalid_rom[  456] = 0; 
    i_addr_rom[  457] = 'h0000004c; 	    d_addr_rom[  457] = 'h00000a40; 	    wdata_rom[  457] = 'hb059c4fa; 	    wvalid_rom[  457] = 0; 
    i_addr_rom[  458] = 'h00000078; 	    d_addr_rom[  458] = 'h00000be4; 	    wdata_rom[  458] = 'h7ed45ebc; 	    wvalid_rom[  458] = 0; 
    i_addr_rom[  459] = 'h00000734; 	    d_addr_rom[  459] = 'h000008b4; 	    wdata_rom[  459] = 'hce6f7ccc; 	    wvalid_rom[  459] = 1; 
    i_addr_rom[  460] = 'h000005b0; 	    d_addr_rom[  460] = 'h00000abc; 	    wdata_rom[  460] = 'h633f006b; 	    wvalid_rom[  460] = 1; 
    i_addr_rom[  461] = 'h00000030; 	    d_addr_rom[  461] = 'h00000b30; 	    wdata_rom[  461] = 'h67e075f8; 	    wvalid_rom[  461] = 1; 
    i_addr_rom[  462] = 'h000002d8; 	    d_addr_rom[  462] = 'h00000cd8; 	    wdata_rom[  462] = 'hadac85ce; 	    wvalid_rom[  462] = 0; 
    i_addr_rom[  463] = 'h00000598; 	    d_addr_rom[  463] = 'h00000990; 	    wdata_rom[  463] = 'h62d70e52; 	    wvalid_rom[  463] = 0; 
    i_addr_rom[  464] = 'h000007a0; 	    d_addr_rom[  464] = 'h00000eb4; 	    wdata_rom[  464] = 'h370e0d32; 	    wvalid_rom[  464] = 1; 
    i_addr_rom[  465] = 'h00000670; 	    d_addr_rom[  465] = 'h00000d84; 	    wdata_rom[  465] = 'h5a611ac9; 	    wvalid_rom[  465] = 0; 
    i_addr_rom[  466] = 'h00000120; 	    d_addr_rom[  466] = 'h00000f2c; 	    wdata_rom[  466] = 'hc67d68eb; 	    wvalid_rom[  466] = 1; 
    i_addr_rom[  467] = 'h000003cc; 	    d_addr_rom[  467] = 'h00000a44; 	    wdata_rom[  467] = 'h6d91fcb2; 	    wvalid_rom[  467] = 1; 
    i_addr_rom[  468] = 'h000007d4; 	    d_addr_rom[  468] = 'h00000b40; 	    wdata_rom[  468] = 'h1cb5e2d3; 	    wvalid_rom[  468] = 0; 
    i_addr_rom[  469] = 'h000006ec; 	    d_addr_rom[  469] = 'h00000bc0; 	    wdata_rom[  469] = 'h1453ff6a; 	    wvalid_rom[  469] = 0; 
    i_addr_rom[  470] = 'h00000584; 	    d_addr_rom[  470] = 'h000009b8; 	    wdata_rom[  470] = 'h161d9413; 	    wvalid_rom[  470] = 1; 
    i_addr_rom[  471] = 'h0000004c; 	    d_addr_rom[  471] = 'h00000f68; 	    wdata_rom[  471] = 'h2735500c; 	    wvalid_rom[  471] = 1; 
    i_addr_rom[  472] = 'h000002e4; 	    d_addr_rom[  472] = 'h00000fe8; 	    wdata_rom[  472] = 'hd1135fbf; 	    wvalid_rom[  472] = 1; 
    i_addr_rom[  473] = 'h000000c4; 	    d_addr_rom[  473] = 'h00000b4c; 	    wdata_rom[  473] = 'hb8462206; 	    wvalid_rom[  473] = 0; 
    i_addr_rom[  474] = 'h000005bc; 	    d_addr_rom[  474] = 'h000008d8; 	    wdata_rom[  474] = 'h6c3f3496; 	    wvalid_rom[  474] = 1; 
    i_addr_rom[  475] = 'h000006c4; 	    d_addr_rom[  475] = 'h00000ef4; 	    wdata_rom[  475] = 'hc34209c6; 	    wvalid_rom[  475] = 0; 
    i_addr_rom[  476] = 'h000004b8; 	    d_addr_rom[  476] = 'h00000e9c; 	    wdata_rom[  476] = 'h31d07c7c; 	    wvalid_rom[  476] = 0; 
    i_addr_rom[  477] = 'h00000004; 	    d_addr_rom[  477] = 'h00000930; 	    wdata_rom[  477] = 'hd8c571fa; 	    wvalid_rom[  477] = 1; 
    i_addr_rom[  478] = 'h00000598; 	    d_addr_rom[  478] = 'h00000b08; 	    wdata_rom[  478] = 'hedf21c6c; 	    wvalid_rom[  478] = 1; 
    i_addr_rom[  479] = 'h0000032c; 	    d_addr_rom[  479] = 'h00000f20; 	    wdata_rom[  479] = 'h575adc77; 	    wvalid_rom[  479] = 1; 
    i_addr_rom[  480] = 'h00000294; 	    d_addr_rom[  480] = 'h00000ba8; 	    wdata_rom[  480] = 'h035ec35a; 	    wvalid_rom[  480] = 1; 
    i_addr_rom[  481] = 'h000006a8; 	    d_addr_rom[  481] = 'h00000e20; 	    wdata_rom[  481] = 'h951d9272; 	    wvalid_rom[  481] = 1; 
    i_addr_rom[  482] = 'h000002e8; 	    d_addr_rom[  482] = 'h00000b0c; 	    wdata_rom[  482] = 'h219bba6f; 	    wvalid_rom[  482] = 0; 
    i_addr_rom[  483] = 'h000004c4; 	    d_addr_rom[  483] = 'h00000bcc; 	    wdata_rom[  483] = 'h1b4272e3; 	    wvalid_rom[  483] = 0; 
    i_addr_rom[  484] = 'h0000041c; 	    d_addr_rom[  484] = 'h00000a38; 	    wdata_rom[  484] = 'h8e53e108; 	    wvalid_rom[  484] = 0; 
    i_addr_rom[  485] = 'h000005ec; 	    d_addr_rom[  485] = 'h00000e9c; 	    wdata_rom[  485] = 'hf4f712ed; 	    wvalid_rom[  485] = 0; 
    i_addr_rom[  486] = 'h00000750; 	    d_addr_rom[  486] = 'h00000864; 	    wdata_rom[  486] = 'hd0d1d413; 	    wvalid_rom[  486] = 1; 
    i_addr_rom[  487] = 'h000003b0; 	    d_addr_rom[  487] = 'h00000c30; 	    wdata_rom[  487] = 'h1d3c18dc; 	    wvalid_rom[  487] = 1; 
    i_addr_rom[  488] = 'h00000280; 	    d_addr_rom[  488] = 'h00000bc8; 	    wdata_rom[  488] = 'h69e50806; 	    wvalid_rom[  488] = 1; 
    i_addr_rom[  489] = 'h0000040c; 	    d_addr_rom[  489] = 'h00000fd4; 	    wdata_rom[  489] = 'hb77b7ae2; 	    wvalid_rom[  489] = 0; 
    i_addr_rom[  490] = 'h000004e8; 	    d_addr_rom[  490] = 'h00000b04; 	    wdata_rom[  490] = 'h0d642f05; 	    wvalid_rom[  490] = 0; 
    i_addr_rom[  491] = 'h00000518; 	    d_addr_rom[  491] = 'h00000ce8; 	    wdata_rom[  491] = 'h0b734964; 	    wvalid_rom[  491] = 0; 
    i_addr_rom[  492] = 'h00000178; 	    d_addr_rom[  492] = 'h00000a48; 	    wdata_rom[  492] = 'hdad56d52; 	    wvalid_rom[  492] = 1; 
    i_addr_rom[  493] = 'h00000384; 	    d_addr_rom[  493] = 'h00000e98; 	    wdata_rom[  493] = 'h319fd45e; 	    wvalid_rom[  493] = 1; 
    i_addr_rom[  494] = 'h00000190; 	    d_addr_rom[  494] = 'h00000890; 	    wdata_rom[  494] = 'h6bc3a93b; 	    wvalid_rom[  494] = 1; 
    i_addr_rom[  495] = 'h00000454; 	    d_addr_rom[  495] = 'h00000ba0; 	    wdata_rom[  495] = 'h7a0ab053; 	    wvalid_rom[  495] = 1; 
    i_addr_rom[  496] = 'h00000400; 	    d_addr_rom[  496] = 'h00000cd4; 	    wdata_rom[  496] = 'hd8f83998; 	    wvalid_rom[  496] = 1; 
    i_addr_rom[  497] = 'h00000170; 	    d_addr_rom[  497] = 'h00000978; 	    wdata_rom[  497] = 'hbe209893; 	    wvalid_rom[  497] = 0; 
    i_addr_rom[  498] = 'h00000254; 	    d_addr_rom[  498] = 'h00000c48; 	    wdata_rom[  498] = 'h00aa246f; 	    wvalid_rom[  498] = 1; 
    i_addr_rom[  499] = 'h00000628; 	    d_addr_rom[  499] = 'h00000ec4; 	    wdata_rom[  499] = 'h93da29a7; 	    wvalid_rom[  499] = 1; 
    i_addr_rom[  500] = 'h00000418; 	    d_addr_rom[  500] = 'h00000820; 	    wdata_rom[  500] = 'h4d8bd26b; 	    wvalid_rom[  500] = 1; 
    i_addr_rom[  501] = 'h00000108; 	    d_addr_rom[  501] = 'h00000ff4; 	    wdata_rom[  501] = 'h15d61bc2; 	    wvalid_rom[  501] = 1; 
    i_addr_rom[  502] = 'h00000028; 	    d_addr_rom[  502] = 'h00000d54; 	    wdata_rom[  502] = 'had319e49; 	    wvalid_rom[  502] = 1; 
    i_addr_rom[  503] = 'h000003c8; 	    d_addr_rom[  503] = 'h00000bc4; 	    wdata_rom[  503] = 'h2c8bc8a4; 	    wvalid_rom[  503] = 0; 
    i_addr_rom[  504] = 'h00000318; 	    d_addr_rom[  504] = 'h00000fe4; 	    wdata_rom[  504] = 'he87a2684; 	    wvalid_rom[  504] = 0; 
    i_addr_rom[  505] = 'h000006d8; 	    d_addr_rom[  505] = 'h00000e14; 	    wdata_rom[  505] = 'hb1974f2c; 	    wvalid_rom[  505] = 0; 
    i_addr_rom[  506] = 'h00000578; 	    d_addr_rom[  506] = 'h00000b4c; 	    wdata_rom[  506] = 'h31619dcd; 	    wvalid_rom[  506] = 1; 
    i_addr_rom[  507] = 'h000006e8; 	    d_addr_rom[  507] = 'h00000a64; 	    wdata_rom[  507] = 'hab5a6e43; 	    wvalid_rom[  507] = 0; 
    i_addr_rom[  508] = 'h00000080; 	    d_addr_rom[  508] = 'h000008c0; 	    wdata_rom[  508] = 'hab20d607; 	    wvalid_rom[  508] = 0; 
    i_addr_rom[  509] = 'h000006bc; 	    d_addr_rom[  509] = 'h00000cf4; 	    wdata_rom[  509] = 'h860cb71c; 	    wvalid_rom[  509] = 0; 
    i_addr_rom[  510] = 'h0000023c; 	    d_addr_rom[  510] = 'h00000c70; 	    wdata_rom[  510] = 'hdc59aa4d; 	    wvalid_rom[  510] = 0; 
    i_addr_rom[  511] = 'h00000310; 	    d_addr_rom[  511] = 'h00000b34; 	    wdata_rom[  511] = 'hc507e858; 	    wvalid_rom[  511] = 1; 
    i_addr_rom[  512] = 'h00000624; 	    d_addr_rom[  512] = 'h00000b2c; 	    wdata_rom[  512] = 'h34dbcad6; 	    wvalid_rom[  512] = 1; 
    i_addr_rom[  513] = 'h000003b4; 	    d_addr_rom[  513] = 'h00000bac; 	    wdata_rom[  513] = 'hc6caad56; 	    wvalid_rom[  513] = 0; 
    i_addr_rom[  514] = 'h00000158; 	    d_addr_rom[  514] = 'h00000f50; 	    wdata_rom[  514] = 'h10b8fd50; 	    wvalid_rom[  514] = 1; 
    i_addr_rom[  515] = 'h000006b8; 	    d_addr_rom[  515] = 'h00000a00; 	    wdata_rom[  515] = 'h8e6aa3e4; 	    wvalid_rom[  515] = 1; 
    i_addr_rom[  516] = 'h000007d4; 	    d_addr_rom[  516] = 'h00000ed8; 	    wdata_rom[  516] = 'h2ff2d6d5; 	    wvalid_rom[  516] = 1; 
    i_addr_rom[  517] = 'h000005e8; 	    d_addr_rom[  517] = 'h00000dd4; 	    wdata_rom[  517] = 'h5d99bdef; 	    wvalid_rom[  517] = 1; 
    i_addr_rom[  518] = 'h000004ec; 	    d_addr_rom[  518] = 'h00000c54; 	    wdata_rom[  518] = 'hbef3dd32; 	    wvalid_rom[  518] = 1; 
    i_addr_rom[  519] = 'h00000728; 	    d_addr_rom[  519] = 'h00000a28; 	    wdata_rom[  519] = 'h2bc20e64; 	    wvalid_rom[  519] = 0; 
    i_addr_rom[  520] = 'h00000488; 	    d_addr_rom[  520] = 'h000008a8; 	    wdata_rom[  520] = 'h97355e96; 	    wvalid_rom[  520] = 1; 
    i_addr_rom[  521] = 'h0000051c; 	    d_addr_rom[  521] = 'h00000abc; 	    wdata_rom[  521] = 'h44502345; 	    wvalid_rom[  521] = 1; 
    i_addr_rom[  522] = 'h000002bc; 	    d_addr_rom[  522] = 'h00000998; 	    wdata_rom[  522] = 'he42a8bd3; 	    wvalid_rom[  522] = 1; 
    i_addr_rom[  523] = 'h000006fc; 	    d_addr_rom[  523] = 'h00000f74; 	    wdata_rom[  523] = 'h9118224a; 	    wvalid_rom[  523] = 1; 
    i_addr_rom[  524] = 'h00000408; 	    d_addr_rom[  524] = 'h00000b24; 	    wdata_rom[  524] = 'hd285f453; 	    wvalid_rom[  524] = 0; 
    i_addr_rom[  525] = 'h000001f8; 	    d_addr_rom[  525] = 'h00000a20; 	    wdata_rom[  525] = 'h0c78d55a; 	    wvalid_rom[  525] = 0; 
    i_addr_rom[  526] = 'h00000094; 	    d_addr_rom[  526] = 'h00000910; 	    wdata_rom[  526] = 'h228994e0; 	    wvalid_rom[  526] = 1; 
    i_addr_rom[  527] = 'h00000738; 	    d_addr_rom[  527] = 'h00000f44; 	    wdata_rom[  527] = 'he0d512c6; 	    wvalid_rom[  527] = 1; 
    i_addr_rom[  528] = 'h00000624; 	    d_addr_rom[  528] = 'h0000089c; 	    wdata_rom[  528] = 'ha5b05e04; 	    wvalid_rom[  528] = 0; 
    i_addr_rom[  529] = 'h000002d8; 	    d_addr_rom[  529] = 'h00000b04; 	    wdata_rom[  529] = 'h33ded1e5; 	    wvalid_rom[  529] = 0; 
    i_addr_rom[  530] = 'h0000021c; 	    d_addr_rom[  530] = 'h000009a4; 	    wdata_rom[  530] = 'h1b1854ee; 	    wvalid_rom[  530] = 1; 
    i_addr_rom[  531] = 'h00000488; 	    d_addr_rom[  531] = 'h0000090c; 	    wdata_rom[  531] = 'h2a58afb8; 	    wvalid_rom[  531] = 0; 
    i_addr_rom[  532] = 'h000003b8; 	    d_addr_rom[  532] = 'h00000d40; 	    wdata_rom[  532] = 'hfb366dd1; 	    wvalid_rom[  532] = 0; 
    i_addr_rom[  533] = 'h000006e0; 	    d_addr_rom[  533] = 'h00000f28; 	    wdata_rom[  533] = 'ha34778ff; 	    wvalid_rom[  533] = 0; 
    i_addr_rom[  534] = 'h00000000; 	    d_addr_rom[  534] = 'h00000b18; 	    wdata_rom[  534] = 'h5c49cbde; 	    wvalid_rom[  534] = 1; 
    i_addr_rom[  535] = 'h000000e4; 	    d_addr_rom[  535] = 'h00000970; 	    wdata_rom[  535] = 'h84ba857b; 	    wvalid_rom[  535] = 0; 
    i_addr_rom[  536] = 'h00000020; 	    d_addr_rom[  536] = 'h00000b40; 	    wdata_rom[  536] = 'hce07c12b; 	    wvalid_rom[  536] = 0; 
    i_addr_rom[  537] = 'h000000f4; 	    d_addr_rom[  537] = 'h00000ca0; 	    wdata_rom[  537] = 'h7ad374d7; 	    wvalid_rom[  537] = 0; 
    i_addr_rom[  538] = 'h000006f8; 	    d_addr_rom[  538] = 'h00000cc8; 	    wdata_rom[  538] = 'heef841fd; 	    wvalid_rom[  538] = 1; 
    i_addr_rom[  539] = 'h00000794; 	    d_addr_rom[  539] = 'h00000988; 	    wdata_rom[  539] = 'he8b2c92d; 	    wvalid_rom[  539] = 1; 
    i_addr_rom[  540] = 'h00000574; 	    d_addr_rom[  540] = 'h00000dfc; 	    wdata_rom[  540] = 'h57560461; 	    wvalid_rom[  540] = 1; 
    i_addr_rom[  541] = 'h0000007c; 	    d_addr_rom[  541] = 'h0000091c; 	    wdata_rom[  541] = 'h165956d8; 	    wvalid_rom[  541] = 0; 
    i_addr_rom[  542] = 'h00000250; 	    d_addr_rom[  542] = 'h00000e9c; 	    wdata_rom[  542] = 'h2f00fb4d; 	    wvalid_rom[  542] = 1; 
    i_addr_rom[  543] = 'h00000548; 	    d_addr_rom[  543] = 'h00000824; 	    wdata_rom[  543] = 'h72a0d2ed; 	    wvalid_rom[  543] = 1; 
    i_addr_rom[  544] = 'h00000574; 	    d_addr_rom[  544] = 'h00000a8c; 	    wdata_rom[  544] = 'h2ce7c229; 	    wvalid_rom[  544] = 1; 
    i_addr_rom[  545] = 'h00000798; 	    d_addr_rom[  545] = 'h00000f30; 	    wdata_rom[  545] = 'h8f9e8c75; 	    wvalid_rom[  545] = 0; 
    i_addr_rom[  546] = 'h000007c8; 	    d_addr_rom[  546] = 'h000008e0; 	    wdata_rom[  546] = 'hc94a5f82; 	    wvalid_rom[  546] = 0; 
    i_addr_rom[  547] = 'h000001e4; 	    d_addr_rom[  547] = 'h00000b84; 	    wdata_rom[  547] = 'hecc7249c; 	    wvalid_rom[  547] = 1; 
    i_addr_rom[  548] = 'h00000038; 	    d_addr_rom[  548] = 'h0000082c; 	    wdata_rom[  548] = 'h17134472; 	    wvalid_rom[  548] = 0; 
    i_addr_rom[  549] = 'h0000031c; 	    d_addr_rom[  549] = 'h00000e14; 	    wdata_rom[  549] = 'h42c5885c; 	    wvalid_rom[  549] = 1; 
    i_addr_rom[  550] = 'h00000600; 	    d_addr_rom[  550] = 'h00000ad0; 	    wdata_rom[  550] = 'h830927f8; 	    wvalid_rom[  550] = 0; 
    i_addr_rom[  551] = 'h00000524; 	    d_addr_rom[  551] = 'h00000a70; 	    wdata_rom[  551] = 'h0257ed29; 	    wvalid_rom[  551] = 0; 
    i_addr_rom[  552] = 'h000003a8; 	    d_addr_rom[  552] = 'h00000b20; 	    wdata_rom[  552] = 'hb210d169; 	    wvalid_rom[  552] = 0; 
    i_addr_rom[  553] = 'h000006f4; 	    d_addr_rom[  553] = 'h00000e40; 	    wdata_rom[  553] = 'h9c7ee0f3; 	    wvalid_rom[  553] = 0; 
    i_addr_rom[  554] = 'h0000067c; 	    d_addr_rom[  554] = 'h00000f64; 	    wdata_rom[  554] = 'hf9024b2c; 	    wvalid_rom[  554] = 1; 
    i_addr_rom[  555] = 'h0000018c; 	    d_addr_rom[  555] = 'h00000ce0; 	    wdata_rom[  555] = 'h3f9ce0a3; 	    wvalid_rom[  555] = 0; 
    i_addr_rom[  556] = 'h000007f0; 	    d_addr_rom[  556] = 'h00000d44; 	    wdata_rom[  556] = 'hcaae4d13; 	    wvalid_rom[  556] = 1; 
    i_addr_rom[  557] = 'h00000538; 	    d_addr_rom[  557] = 'h00000ecc; 	    wdata_rom[  557] = 'h241f0f9b; 	    wvalid_rom[  557] = 0; 
    i_addr_rom[  558] = 'h000006f8; 	    d_addr_rom[  558] = 'h00000bac; 	    wdata_rom[  558] = 'haff07706; 	    wvalid_rom[  558] = 0; 
    i_addr_rom[  559] = 'h00000034; 	    d_addr_rom[  559] = 'h00000e0c; 	    wdata_rom[  559] = 'h6c15a766; 	    wvalid_rom[  559] = 1; 
    i_addr_rom[  560] = 'h0000046c; 	    d_addr_rom[  560] = 'h00000a14; 	    wdata_rom[  560] = 'h7c131ad8; 	    wvalid_rom[  560] = 0; 
    i_addr_rom[  561] = 'h0000060c; 	    d_addr_rom[  561] = 'h0000086c; 	    wdata_rom[  561] = 'h4713ac94; 	    wvalid_rom[  561] = 0; 
    i_addr_rom[  562] = 'h000002d8; 	    d_addr_rom[  562] = 'h00000904; 	    wdata_rom[  562] = 'h7f2d75a6; 	    wvalid_rom[  562] = 0; 
    i_addr_rom[  563] = 'h00000604; 	    d_addr_rom[  563] = 'h00000a04; 	    wdata_rom[  563] = 'h3df49b61; 	    wvalid_rom[  563] = 0; 
    i_addr_rom[  564] = 'h0000008c; 	    d_addr_rom[  564] = 'h00000b84; 	    wdata_rom[  564] = 'hf76aa257; 	    wvalid_rom[  564] = 0; 
    i_addr_rom[  565] = 'h00000134; 	    d_addr_rom[  565] = 'h00000d1c; 	    wdata_rom[  565] = 'h89130a25; 	    wvalid_rom[  565] = 1; 
    i_addr_rom[  566] = 'h000006d4; 	    d_addr_rom[  566] = 'h00000fa8; 	    wdata_rom[  566] = 'ha13172cb; 	    wvalid_rom[  566] = 0; 
    i_addr_rom[  567] = 'h000001d4; 	    d_addr_rom[  567] = 'h00000cd4; 	    wdata_rom[  567] = 'h41d0c653; 	    wvalid_rom[  567] = 1; 
    i_addr_rom[  568] = 'h00000690; 	    d_addr_rom[  568] = 'h00000c54; 	    wdata_rom[  568] = 'h66831d35; 	    wvalid_rom[  568] = 1; 
    i_addr_rom[  569] = 'h00000210; 	    d_addr_rom[  569] = 'h00000e98; 	    wdata_rom[  569] = 'hc6fcca15; 	    wvalid_rom[  569] = 0; 
    i_addr_rom[  570] = 'h00000380; 	    d_addr_rom[  570] = 'h00000aa0; 	    wdata_rom[  570] = 'h9d165b2c; 	    wvalid_rom[  570] = 0; 
    i_addr_rom[  571] = 'h000007a8; 	    d_addr_rom[  571] = 'h00000a40; 	    wdata_rom[  571] = 'h1a36879e; 	    wvalid_rom[  571] = 1; 
    i_addr_rom[  572] = 'h00000354; 	    d_addr_rom[  572] = 'h000008f8; 	    wdata_rom[  572] = 'h541c462e; 	    wvalid_rom[  572] = 0; 
    i_addr_rom[  573] = 'h000003a0; 	    d_addr_rom[  573] = 'h00000fe4; 	    wdata_rom[  573] = 'h20666cb6; 	    wvalid_rom[  573] = 1; 
    i_addr_rom[  574] = 'h00000614; 	    d_addr_rom[  574] = 'h00000860; 	    wdata_rom[  574] = 'h4abd6d7f; 	    wvalid_rom[  574] = 0; 
    i_addr_rom[  575] = 'h00000074; 	    d_addr_rom[  575] = 'h000009fc; 	    wdata_rom[  575] = 'h76bf9c7f; 	    wvalid_rom[  575] = 0; 
    i_addr_rom[  576] = 'h0000050c; 	    d_addr_rom[  576] = 'h00000e2c; 	    wdata_rom[  576] = 'hda52dc2a; 	    wvalid_rom[  576] = 1; 
    i_addr_rom[  577] = 'h00000220; 	    d_addr_rom[  577] = 'h0000084c; 	    wdata_rom[  577] = 'h78504c88; 	    wvalid_rom[  577] = 1; 
    i_addr_rom[  578] = 'h000004d4; 	    d_addr_rom[  578] = 'h00000d64; 	    wdata_rom[  578] = 'hbfe580d2; 	    wvalid_rom[  578] = 0; 
    i_addr_rom[  579] = 'h0000029c; 	    d_addr_rom[  579] = 'h00000fcc; 	    wdata_rom[  579] = 'hd3dc2531; 	    wvalid_rom[  579] = 1; 
    i_addr_rom[  580] = 'h0000035c; 	    d_addr_rom[  580] = 'h00000c3c; 	    wdata_rom[  580] = 'h96a25f68; 	    wvalid_rom[  580] = 1; 
    i_addr_rom[  581] = 'h000006c4; 	    d_addr_rom[  581] = 'h00000a8c; 	    wdata_rom[  581] = 'h32d388da; 	    wvalid_rom[  581] = 0; 
    i_addr_rom[  582] = 'h0000068c; 	    d_addr_rom[  582] = 'h00000a4c; 	    wdata_rom[  582] = 'hcf54dc85; 	    wvalid_rom[  582] = 0; 
    i_addr_rom[  583] = 'h0000030c; 	    d_addr_rom[  583] = 'h00000ce8; 	    wdata_rom[  583] = 'h06e78084; 	    wvalid_rom[  583] = 1; 
    i_addr_rom[  584] = 'h000003d0; 	    d_addr_rom[  584] = 'h00000f84; 	    wdata_rom[  584] = 'h168d7d8f; 	    wvalid_rom[  584] = 1; 
    i_addr_rom[  585] = 'h000007b4; 	    d_addr_rom[  585] = 'h0000085c; 	    wdata_rom[  585] = 'h7d0c8553; 	    wvalid_rom[  585] = 1; 
    i_addr_rom[  586] = 'h000002c0; 	    d_addr_rom[  586] = 'h00000d70; 	    wdata_rom[  586] = 'hde2f56e9; 	    wvalid_rom[  586] = 0; 
    i_addr_rom[  587] = 'h00000114; 	    d_addr_rom[  587] = 'h00000f40; 	    wdata_rom[  587] = 'hee3e826f; 	    wvalid_rom[  587] = 1; 
    i_addr_rom[  588] = 'h0000029c; 	    d_addr_rom[  588] = 'h00000cd4; 	    wdata_rom[  588] = 'h03b5d948; 	    wvalid_rom[  588] = 0; 
    i_addr_rom[  589] = 'h000001d0; 	    d_addr_rom[  589] = 'h00000c48; 	    wdata_rom[  589] = 'he22c1f75; 	    wvalid_rom[  589] = 1; 
    i_addr_rom[  590] = 'h00000780; 	    d_addr_rom[  590] = 'h00000ab8; 	    wdata_rom[  590] = 'h4b3f5a77; 	    wvalid_rom[  590] = 1; 
    i_addr_rom[  591] = 'h000005d4; 	    d_addr_rom[  591] = 'h00000f54; 	    wdata_rom[  591] = 'h45c6e922; 	    wvalid_rom[  591] = 0; 
    i_addr_rom[  592] = 'h00000568; 	    d_addr_rom[  592] = 'h00000f88; 	    wdata_rom[  592] = 'h839d2399; 	    wvalid_rom[  592] = 0; 
    i_addr_rom[  593] = 'h000005ec; 	    d_addr_rom[  593] = 'h00000a7c; 	    wdata_rom[  593] = 'h2606a0a2; 	    wvalid_rom[  593] = 0; 
    i_addr_rom[  594] = 'h000005d4; 	    d_addr_rom[  594] = 'h00000f0c; 	    wdata_rom[  594] = 'haccac797; 	    wvalid_rom[  594] = 1; 
    i_addr_rom[  595] = 'h0000071c; 	    d_addr_rom[  595] = 'h00000d00; 	    wdata_rom[  595] = 'h6ac15b99; 	    wvalid_rom[  595] = 1; 
    i_addr_rom[  596] = 'h00000458; 	    d_addr_rom[  596] = 'h000008f8; 	    wdata_rom[  596] = 'he7076f53; 	    wvalid_rom[  596] = 1; 
    i_addr_rom[  597] = 'h00000360; 	    d_addr_rom[  597] = 'h00000d04; 	    wdata_rom[  597] = 'h21a53280; 	    wvalid_rom[  597] = 0; 
    i_addr_rom[  598] = 'h000007bc; 	    d_addr_rom[  598] = 'h000009bc; 	    wdata_rom[  598] = 'haa917a53; 	    wvalid_rom[  598] = 1; 
    i_addr_rom[  599] = 'h000005fc; 	    d_addr_rom[  599] = 'h00000e64; 	    wdata_rom[  599] = 'h1bcf8d92; 	    wvalid_rom[  599] = 0; 
    i_addr_rom[  600] = 'h0000065c; 	    d_addr_rom[  600] = 'h00000d78; 	    wdata_rom[  600] = 'h8ea6ce25; 	    wvalid_rom[  600] = 1; 
    i_addr_rom[  601] = 'h00000700; 	    d_addr_rom[  601] = 'h00000838; 	    wdata_rom[  601] = 'hb66052e5; 	    wvalid_rom[  601] = 1; 
    i_addr_rom[  602] = 'h00000024; 	    d_addr_rom[  602] = 'h00000b48; 	    wdata_rom[  602] = 'h51da4c1f; 	    wvalid_rom[  602] = 0; 
    i_addr_rom[  603] = 'h000006ac; 	    d_addr_rom[  603] = 'h00000c28; 	    wdata_rom[  603] = 'h24260e0b; 	    wvalid_rom[  603] = 0; 
    i_addr_rom[  604] = 'h0000059c; 	    d_addr_rom[  604] = 'h00000bd0; 	    wdata_rom[  604] = 'he1f509a5; 	    wvalid_rom[  604] = 0; 
    i_addr_rom[  605] = 'h000004ec; 	    d_addr_rom[  605] = 'h00000870; 	    wdata_rom[  605] = 'hdc6f62ac; 	    wvalid_rom[  605] = 1; 
    i_addr_rom[  606] = 'h0000067c; 	    d_addr_rom[  606] = 'h00000ed0; 	    wdata_rom[  606] = 'h10b918b3; 	    wvalid_rom[  606] = 0; 
    i_addr_rom[  607] = 'h0000021c; 	    d_addr_rom[  607] = 'h00000f10; 	    wdata_rom[  607] = 'he2bce631; 	    wvalid_rom[  607] = 0; 
    i_addr_rom[  608] = 'h00000218; 	    d_addr_rom[  608] = 'h00000844; 	    wdata_rom[  608] = 'he4113a6a; 	    wvalid_rom[  608] = 1; 
    i_addr_rom[  609] = 'h00000610; 	    d_addr_rom[  609] = 'h00000918; 	    wdata_rom[  609] = 'h0f2b5bf7; 	    wvalid_rom[  609] = 0; 
    i_addr_rom[  610] = 'h00000394; 	    d_addr_rom[  610] = 'h00000d0c; 	    wdata_rom[  610] = 'h6e77cd0d; 	    wvalid_rom[  610] = 1; 
    i_addr_rom[  611] = 'h000004f4; 	    d_addr_rom[  611] = 'h0000091c; 	    wdata_rom[  611] = 'h185a1397; 	    wvalid_rom[  611] = 0; 
    i_addr_rom[  612] = 'h0000028c; 	    d_addr_rom[  612] = 'h00000ee8; 	    wdata_rom[  612] = 'hf295a446; 	    wvalid_rom[  612] = 0; 
    i_addr_rom[  613] = 'h00000408; 	    d_addr_rom[  613] = 'h00000c24; 	    wdata_rom[  613] = 'hbc4bd17a; 	    wvalid_rom[  613] = 0; 
    i_addr_rom[  614] = 'h00000690; 	    d_addr_rom[  614] = 'h00000f88; 	    wdata_rom[  614] = 'hecd6f149; 	    wvalid_rom[  614] = 0; 
    i_addr_rom[  615] = 'h00000494; 	    d_addr_rom[  615] = 'h00000c80; 	    wdata_rom[  615] = 'h52b2649c; 	    wvalid_rom[  615] = 1; 
    i_addr_rom[  616] = 'h00000794; 	    d_addr_rom[  616] = 'h00000bcc; 	    wdata_rom[  616] = 'hc56c3330; 	    wvalid_rom[  616] = 0; 
    i_addr_rom[  617] = 'h00000388; 	    d_addr_rom[  617] = 'h00000e14; 	    wdata_rom[  617] = 'h0ac005ed; 	    wvalid_rom[  617] = 1; 
    i_addr_rom[  618] = 'h00000138; 	    d_addr_rom[  618] = 'h000009dc; 	    wdata_rom[  618] = 'h1286e9a2; 	    wvalid_rom[  618] = 0; 
    i_addr_rom[  619] = 'h00000564; 	    d_addr_rom[  619] = 'h00000830; 	    wdata_rom[  619] = 'hfdf6ee56; 	    wvalid_rom[  619] = 0; 
    i_addr_rom[  620] = 'h00000174; 	    d_addr_rom[  620] = 'h00000b2c; 	    wdata_rom[  620] = 'h8b1551e6; 	    wvalid_rom[  620] = 1; 
    i_addr_rom[  621] = 'h0000027c; 	    d_addr_rom[  621] = 'h00000c2c; 	    wdata_rom[  621] = 'h06684585; 	    wvalid_rom[  621] = 1; 
    i_addr_rom[  622] = 'h00000600; 	    d_addr_rom[  622] = 'h00000d54; 	    wdata_rom[  622] = 'h1e7416d2; 	    wvalid_rom[  622] = 0; 
    i_addr_rom[  623] = 'h000004d0; 	    d_addr_rom[  623] = 'h00000dd8; 	    wdata_rom[  623] = 'h4a067858; 	    wvalid_rom[  623] = 0; 
    i_addr_rom[  624] = 'h000007d0; 	    d_addr_rom[  624] = 'h00000d68; 	    wdata_rom[  624] = 'h84da2def; 	    wvalid_rom[  624] = 0; 
    i_addr_rom[  625] = 'h00000154; 	    d_addr_rom[  625] = 'h00000974; 	    wdata_rom[  625] = 'hfb4f8f19; 	    wvalid_rom[  625] = 1; 
    i_addr_rom[  626] = 'h00000330; 	    d_addr_rom[  626] = 'h00000d4c; 	    wdata_rom[  626] = 'haffa5bdc; 	    wvalid_rom[  626] = 0; 
    i_addr_rom[  627] = 'h0000059c; 	    d_addr_rom[  627] = 'h000008e8; 	    wdata_rom[  627] = 'h340c77ca; 	    wvalid_rom[  627] = 1; 
    i_addr_rom[  628] = 'h00000168; 	    d_addr_rom[  628] = 'h000009e0; 	    wdata_rom[  628] = 'hc86efe62; 	    wvalid_rom[  628] = 0; 
    i_addr_rom[  629] = 'h000004a0; 	    d_addr_rom[  629] = 'h00000c64; 	    wdata_rom[  629] = 'h6b8e990f; 	    wvalid_rom[  629] = 0; 
    i_addr_rom[  630] = 'h000001f8; 	    d_addr_rom[  630] = 'h00000c40; 	    wdata_rom[  630] = 'h2a4589c4; 	    wvalid_rom[  630] = 0; 
    i_addr_rom[  631] = 'h000002fc; 	    d_addr_rom[  631] = 'h000008cc; 	    wdata_rom[  631] = 'hb311727e; 	    wvalid_rom[  631] = 0; 
    i_addr_rom[  632] = 'h000007b0; 	    d_addr_rom[  632] = 'h00000e74; 	    wdata_rom[  632] = 'h5ed59530; 	    wvalid_rom[  632] = 1; 
    i_addr_rom[  633] = 'h00000128; 	    d_addr_rom[  633] = 'h00000a04; 	    wdata_rom[  633] = 'he3bce97b; 	    wvalid_rom[  633] = 0; 
    i_addr_rom[  634] = 'h000000b4; 	    d_addr_rom[  634] = 'h00000890; 	    wdata_rom[  634] = 'hb2135e32; 	    wvalid_rom[  634] = 0; 
    i_addr_rom[  635] = 'h00000394; 	    d_addr_rom[  635] = 'h00000ecc; 	    wdata_rom[  635] = 'h36404e3b; 	    wvalid_rom[  635] = 0; 
    i_addr_rom[  636] = 'h00000310; 	    d_addr_rom[  636] = 'h00000ef0; 	    wdata_rom[  636] = 'hf6956307; 	    wvalid_rom[  636] = 0; 
    i_addr_rom[  637] = 'h00000114; 	    d_addr_rom[  637] = 'h00000820; 	    wdata_rom[  637] = 'hf8ef2bfa; 	    wvalid_rom[  637] = 0; 
    i_addr_rom[  638] = 'h00000074; 	    d_addr_rom[  638] = 'h00000e1c; 	    wdata_rom[  638] = 'h8c21723e; 	    wvalid_rom[  638] = 1; 
    i_addr_rom[  639] = 'h00000700; 	    d_addr_rom[  639] = 'h00000bc8; 	    wdata_rom[  639] = 'h976c2167; 	    wvalid_rom[  639] = 1; 
    i_addr_rom[  640] = 'h00000554; 	    d_addr_rom[  640] = 'h00000f20; 	    wdata_rom[  640] = 'hc5de785d; 	    wvalid_rom[  640] = 1; 
    i_addr_rom[  641] = 'h0000004c; 	    d_addr_rom[  641] = 'h00000de0; 	    wdata_rom[  641] = 'hdaca4f49; 	    wvalid_rom[  641] = 0; 
    i_addr_rom[  642] = 'h00000214; 	    d_addr_rom[  642] = 'h00000b10; 	    wdata_rom[  642] = 'ha06aa68e; 	    wvalid_rom[  642] = 1; 
    i_addr_rom[  643] = 'h000006c8; 	    d_addr_rom[  643] = 'h00000a88; 	    wdata_rom[  643] = 'h8bd13286; 	    wvalid_rom[  643] = 0; 
    i_addr_rom[  644] = 'h0000005c; 	    d_addr_rom[  644] = 'h00000bd8; 	    wdata_rom[  644] = 'h529de99a; 	    wvalid_rom[  644] = 1; 
    i_addr_rom[  645] = 'h00000170; 	    d_addr_rom[  645] = 'h00000ba8; 	    wdata_rom[  645] = 'h098b9d32; 	    wvalid_rom[  645] = 1; 
    i_addr_rom[  646] = 'h00000670; 	    d_addr_rom[  646] = 'h00000d70; 	    wdata_rom[  646] = 'h8c3a3e53; 	    wvalid_rom[  646] = 0; 
    i_addr_rom[  647] = 'h000000a0; 	    d_addr_rom[  647] = 'h00000b54; 	    wdata_rom[  647] = 'h47bbc93b; 	    wvalid_rom[  647] = 0; 
    i_addr_rom[  648] = 'h00000474; 	    d_addr_rom[  648] = 'h00000b50; 	    wdata_rom[  648] = 'h91f36825; 	    wvalid_rom[  648] = 0; 
    i_addr_rom[  649] = 'h00000644; 	    d_addr_rom[  649] = 'h00000a1c; 	    wdata_rom[  649] = 'h8556c681; 	    wvalid_rom[  649] = 1; 
    i_addr_rom[  650] = 'h000006f4; 	    d_addr_rom[  650] = 'h00000e20; 	    wdata_rom[  650] = 'hab4a189c; 	    wvalid_rom[  650] = 1; 
    i_addr_rom[  651] = 'h000002a4; 	    d_addr_rom[  651] = 'h000009cc; 	    wdata_rom[  651] = 'ha56fa39a; 	    wvalid_rom[  651] = 1; 
    i_addr_rom[  652] = 'h000007f8; 	    d_addr_rom[  652] = 'h00000c64; 	    wdata_rom[  652] = 'h270cd5a3; 	    wvalid_rom[  652] = 0; 
    i_addr_rom[  653] = 'h0000002c; 	    d_addr_rom[  653] = 'h00000de4; 	    wdata_rom[  653] = 'hcfc86e17; 	    wvalid_rom[  653] = 0; 
    i_addr_rom[  654] = 'h000002b4; 	    d_addr_rom[  654] = 'h00000a8c; 	    wdata_rom[  654] = 'h67232919; 	    wvalid_rom[  654] = 1; 
    i_addr_rom[  655] = 'h00000320; 	    d_addr_rom[  655] = 'h00000ab0; 	    wdata_rom[  655] = 'h94ac820b; 	    wvalid_rom[  655] = 1; 
    i_addr_rom[  656] = 'h0000059c; 	    d_addr_rom[  656] = 'h00000b34; 	    wdata_rom[  656] = 'hda835016; 	    wvalid_rom[  656] = 0; 
    i_addr_rom[  657] = 'h000004e0; 	    d_addr_rom[  657] = 'h00000b40; 	    wdata_rom[  657] = 'h39aa173e; 	    wvalid_rom[  657] = 0; 
    i_addr_rom[  658] = 'h0000041c; 	    d_addr_rom[  658] = 'h00000fb0; 	    wdata_rom[  658] = 'h4eff8712; 	    wvalid_rom[  658] = 0; 
    i_addr_rom[  659] = 'h00000360; 	    d_addr_rom[  659] = 'h00000d28; 	    wdata_rom[  659] = 'h50722ec7; 	    wvalid_rom[  659] = 0; 
    i_addr_rom[  660] = 'h00000690; 	    d_addr_rom[  660] = 'h00000c70; 	    wdata_rom[  660] = 'hc85615fe; 	    wvalid_rom[  660] = 1; 
    i_addr_rom[  661] = 'h00000224; 	    d_addr_rom[  661] = 'h00000ca8; 	    wdata_rom[  661] = 'h25794e48; 	    wvalid_rom[  661] = 1; 
    i_addr_rom[  662] = 'h0000001c; 	    d_addr_rom[  662] = 'h000009dc; 	    wdata_rom[  662] = 'h3db3ef79; 	    wvalid_rom[  662] = 1; 
    i_addr_rom[  663] = 'h00000144; 	    d_addr_rom[  663] = 'h00000bd8; 	    wdata_rom[  663] = 'h8ebe4e53; 	    wvalid_rom[  663] = 0; 
    i_addr_rom[  664] = 'h00000234; 	    d_addr_rom[  664] = 'h00000ad8; 	    wdata_rom[  664] = 'h9d170ac3; 	    wvalid_rom[  664] = 1; 
    i_addr_rom[  665] = 'h000001a8; 	    d_addr_rom[  665] = 'h00000a48; 	    wdata_rom[  665] = 'he00e5467; 	    wvalid_rom[  665] = 0; 
    i_addr_rom[  666] = 'h00000178; 	    d_addr_rom[  666] = 'h00000d1c; 	    wdata_rom[  666] = 'hedabdd8d; 	    wvalid_rom[  666] = 0; 
    i_addr_rom[  667] = 'h00000230; 	    d_addr_rom[  667] = 'h00000f7c; 	    wdata_rom[  667] = 'h56505709; 	    wvalid_rom[  667] = 1; 
    i_addr_rom[  668] = 'h000000ac; 	    d_addr_rom[  668] = 'h00000a78; 	    wdata_rom[  668] = 'h1b3ed992; 	    wvalid_rom[  668] = 1; 
    i_addr_rom[  669] = 'h000001d8; 	    d_addr_rom[  669] = 'h00000fe4; 	    wdata_rom[  669] = 'h507f2149; 	    wvalid_rom[  669] = 1; 
    i_addr_rom[  670] = 'h00000150; 	    d_addr_rom[  670] = 'h00000b88; 	    wdata_rom[  670] = 'h2fed7940; 	    wvalid_rom[  670] = 1; 
    i_addr_rom[  671] = 'h000003e0; 	    d_addr_rom[  671] = 'h00000fac; 	    wdata_rom[  671] = 'h91c1746e; 	    wvalid_rom[  671] = 1; 
    i_addr_rom[  672] = 'h000002d0; 	    d_addr_rom[  672] = 'h00000b78; 	    wdata_rom[  672] = 'hb101a280; 	    wvalid_rom[  672] = 1; 
    i_addr_rom[  673] = 'h0000049c; 	    d_addr_rom[  673] = 'h00000bbc; 	    wdata_rom[  673] = 'hce1e004d; 	    wvalid_rom[  673] = 0; 
    i_addr_rom[  674] = 'h00000160; 	    d_addr_rom[  674] = 'h00000e68; 	    wdata_rom[  674] = 'ha2923c92; 	    wvalid_rom[  674] = 1; 
    i_addr_rom[  675] = 'h000001b4; 	    d_addr_rom[  675] = 'h00000830; 	    wdata_rom[  675] = 'h49adcb81; 	    wvalid_rom[  675] = 0; 
    i_addr_rom[  676] = 'h000006b4; 	    d_addr_rom[  676] = 'h00000d74; 	    wdata_rom[  676] = 'h0cba51d2; 	    wvalid_rom[  676] = 1; 
    i_addr_rom[  677] = 'h000007e8; 	    d_addr_rom[  677] = 'h00000d70; 	    wdata_rom[  677] = 'h6099c61f; 	    wvalid_rom[  677] = 1; 
    i_addr_rom[  678] = 'h00000428; 	    d_addr_rom[  678] = 'h00000818; 	    wdata_rom[  678] = 'hf36993d3; 	    wvalid_rom[  678] = 1; 
    i_addr_rom[  679] = 'h0000033c; 	    d_addr_rom[  679] = 'h00000ef0; 	    wdata_rom[  679] = 'h2c1f51f3; 	    wvalid_rom[  679] = 1; 
    i_addr_rom[  680] = 'h0000034c; 	    d_addr_rom[  680] = 'h00000af8; 	    wdata_rom[  680] = 'h6f09d4f3; 	    wvalid_rom[  680] = 0; 
    i_addr_rom[  681] = 'h000001a0; 	    d_addr_rom[  681] = 'h00000ccc; 	    wdata_rom[  681] = 'habfe09b1; 	    wvalid_rom[  681] = 0; 
    i_addr_rom[  682] = 'h00000474; 	    d_addr_rom[  682] = 'h00000d90; 	    wdata_rom[  682] = 'h1343c349; 	    wvalid_rom[  682] = 0; 
    i_addr_rom[  683] = 'h00000008; 	    d_addr_rom[  683] = 'h00000d40; 	    wdata_rom[  683] = 'h0d39ff31; 	    wvalid_rom[  683] = 1; 
    i_addr_rom[  684] = 'h000003a4; 	    d_addr_rom[  684] = 'h00000fe0; 	    wdata_rom[  684] = 'hf820d486; 	    wvalid_rom[  684] = 1; 
    i_addr_rom[  685] = 'h0000059c; 	    d_addr_rom[  685] = 'h00000a80; 	    wdata_rom[  685] = 'ha3fde64c; 	    wvalid_rom[  685] = 0; 
    i_addr_rom[  686] = 'h00000050; 	    d_addr_rom[  686] = 'h00000fd8; 	    wdata_rom[  686] = 'h4aae7387; 	    wvalid_rom[  686] = 0; 
    i_addr_rom[  687] = 'h00000264; 	    d_addr_rom[  687] = 'h00000f58; 	    wdata_rom[  687] = 'hf9f8ab12; 	    wvalid_rom[  687] = 1; 
    i_addr_rom[  688] = 'h000002c4; 	    d_addr_rom[  688] = 'h000008a8; 	    wdata_rom[  688] = 'h2dd37f91; 	    wvalid_rom[  688] = 0; 
    i_addr_rom[  689] = 'h00000790; 	    d_addr_rom[  689] = 'h00000d60; 	    wdata_rom[  689] = 'hcfd63a13; 	    wvalid_rom[  689] = 0; 
    i_addr_rom[  690] = 'h000002a0; 	    d_addr_rom[  690] = 'h00000a74; 	    wdata_rom[  690] = 'hfd44246d; 	    wvalid_rom[  690] = 1; 
    i_addr_rom[  691] = 'h0000032c; 	    d_addr_rom[  691] = 'h000009e4; 	    wdata_rom[  691] = 'heea40893; 	    wvalid_rom[  691] = 1; 
    i_addr_rom[  692] = 'h00000138; 	    d_addr_rom[  692] = 'h00000864; 	    wdata_rom[  692] = 'h0b6e9a11; 	    wvalid_rom[  692] = 0; 
    i_addr_rom[  693] = 'h000006e8; 	    d_addr_rom[  693] = 'h00000e4c; 	    wdata_rom[  693] = 'h3a4a6656; 	    wvalid_rom[  693] = 0; 
    i_addr_rom[  694] = 'h00000610; 	    d_addr_rom[  694] = 'h00000a10; 	    wdata_rom[  694] = 'hd64e8771; 	    wvalid_rom[  694] = 0; 
    i_addr_rom[  695] = 'h00000424; 	    d_addr_rom[  695] = 'h00000efc; 	    wdata_rom[  695] = 'h871ba40c; 	    wvalid_rom[  695] = 1; 
    i_addr_rom[  696] = 'h000003c0; 	    d_addr_rom[  696] = 'h00000840; 	    wdata_rom[  696] = 'hf9d45d01; 	    wvalid_rom[  696] = 0; 
    i_addr_rom[  697] = 'h00000784; 	    d_addr_rom[  697] = 'h00000a20; 	    wdata_rom[  697] = 'h2dcdb8f2; 	    wvalid_rom[  697] = 1; 
    i_addr_rom[  698] = 'h000000d4; 	    d_addr_rom[  698] = 'h00000dec; 	    wdata_rom[  698] = 'h3132610a; 	    wvalid_rom[  698] = 0; 
    i_addr_rom[  699] = 'h000000dc; 	    d_addr_rom[  699] = 'h00000aa0; 	    wdata_rom[  699] = 'h43dace6d; 	    wvalid_rom[  699] = 0; 
    i_addr_rom[  700] = 'h000007e8; 	    d_addr_rom[  700] = 'h00000ed0; 	    wdata_rom[  700] = 'hb2d38ebb; 	    wvalid_rom[  700] = 0; 
    i_addr_rom[  701] = 'h000004a8; 	    d_addr_rom[  701] = 'h00000c9c; 	    wdata_rom[  701] = 'h0af2a3e3; 	    wvalid_rom[  701] = 0; 
    i_addr_rom[  702] = 'h000004e4; 	    d_addr_rom[  702] = 'h000008a0; 	    wdata_rom[  702] = 'h7422f27b; 	    wvalid_rom[  702] = 1; 
    i_addr_rom[  703] = 'h00000424; 	    d_addr_rom[  703] = 'h00000bfc; 	    wdata_rom[  703] = 'hbce15ceb; 	    wvalid_rom[  703] = 0; 
    i_addr_rom[  704] = 'h00000278; 	    d_addr_rom[  704] = 'h00000eec; 	    wdata_rom[  704] = 'he0410caa; 	    wvalid_rom[  704] = 0; 
    i_addr_rom[  705] = 'h0000050c; 	    d_addr_rom[  705] = 'h00000c94; 	    wdata_rom[  705] = 'h91ef1027; 	    wvalid_rom[  705] = 1; 
    i_addr_rom[  706] = 'h00000178; 	    d_addr_rom[  706] = 'h00000a90; 	    wdata_rom[  706] = 'h19c520e6; 	    wvalid_rom[  706] = 0; 
    i_addr_rom[  707] = 'h0000057c; 	    d_addr_rom[  707] = 'h00000e68; 	    wdata_rom[  707] = 'ha292ca1f; 	    wvalid_rom[  707] = 1; 
    i_addr_rom[  708] = 'h000004c0; 	    d_addr_rom[  708] = 'h00000a10; 	    wdata_rom[  708] = 'h6a555854; 	    wvalid_rom[  708] = 1; 
    i_addr_rom[  709] = 'h000006c0; 	    d_addr_rom[  709] = 'h00000f40; 	    wdata_rom[  709] = 'h4159123a; 	    wvalid_rom[  709] = 0; 
    i_addr_rom[  710] = 'h000006a0; 	    d_addr_rom[  710] = 'h00000bd4; 	    wdata_rom[  710] = 'h9d793553; 	    wvalid_rom[  710] = 0; 
    i_addr_rom[  711] = 'h00000340; 	    d_addr_rom[  711] = 'h00000a60; 	    wdata_rom[  711] = 'heb93656b; 	    wvalid_rom[  711] = 0; 
    i_addr_rom[  712] = 'h00000794; 	    d_addr_rom[  712] = 'h00000d84; 	    wdata_rom[  712] = 'h3c6c16fd; 	    wvalid_rom[  712] = 0; 
    i_addr_rom[  713] = 'h000007a8; 	    d_addr_rom[  713] = 'h00000e38; 	    wdata_rom[  713] = 'h98be631c; 	    wvalid_rom[  713] = 0; 
    i_addr_rom[  714] = 'h000002d0; 	    d_addr_rom[  714] = 'h000009dc; 	    wdata_rom[  714] = 'h4e80452f; 	    wvalid_rom[  714] = 1; 
    i_addr_rom[  715] = 'h0000070c; 	    d_addr_rom[  715] = 'h00000e28; 	    wdata_rom[  715] = 'hb112efe1; 	    wvalid_rom[  715] = 1; 
    i_addr_rom[  716] = 'h000000e8; 	    d_addr_rom[  716] = 'h00000f70; 	    wdata_rom[  716] = 'h3b36a8d4; 	    wvalid_rom[  716] = 1; 
    i_addr_rom[  717] = 'h00000594; 	    d_addr_rom[  717] = 'h00000834; 	    wdata_rom[  717] = 'h7b239043; 	    wvalid_rom[  717] = 0; 
    i_addr_rom[  718] = 'h00000204; 	    d_addr_rom[  718] = 'h00000bb8; 	    wdata_rom[  718] = 'he30dfb1f; 	    wvalid_rom[  718] = 0; 
    i_addr_rom[  719] = 'h000000d0; 	    d_addr_rom[  719] = 'h00000b68; 	    wdata_rom[  719] = 'hada9ad72; 	    wvalid_rom[  719] = 1; 
    i_addr_rom[  720] = 'h00000130; 	    d_addr_rom[  720] = 'h00000a1c; 	    wdata_rom[  720] = 'h2fa62c8e; 	    wvalid_rom[  720] = 1; 
    i_addr_rom[  721] = 'h0000022c; 	    d_addr_rom[  721] = 'h00000a28; 	    wdata_rom[  721] = 'hda9a5206; 	    wvalid_rom[  721] = 1; 
    i_addr_rom[  722] = 'h000000a0; 	    d_addr_rom[  722] = 'h000008c0; 	    wdata_rom[  722] = 'h69133801; 	    wvalid_rom[  722] = 1; 
    i_addr_rom[  723] = 'h00000774; 	    d_addr_rom[  723] = 'h00000998; 	    wdata_rom[  723] = 'h803dbf97; 	    wvalid_rom[  723] = 0; 
    i_addr_rom[  724] = 'h00000004; 	    d_addr_rom[  724] = 'h00000fb8; 	    wdata_rom[  724] = 'hed76470f; 	    wvalid_rom[  724] = 1; 
    i_addr_rom[  725] = 'h00000198; 	    d_addr_rom[  725] = 'h00000c2c; 	    wdata_rom[  725] = 'hef3df437; 	    wvalid_rom[  725] = 0; 
    i_addr_rom[  726] = 'h00000328; 	    d_addr_rom[  726] = 'h00000fe0; 	    wdata_rom[  726] = 'h37223ad8; 	    wvalid_rom[  726] = 1; 
    i_addr_rom[  727] = 'h00000688; 	    d_addr_rom[  727] = 'h00000dcc; 	    wdata_rom[  727] = 'h71fddf6c; 	    wvalid_rom[  727] = 0; 
    i_addr_rom[  728] = 'h000002dc; 	    d_addr_rom[  728] = 'h00000ec8; 	    wdata_rom[  728] = 'hbedbaa03; 	    wvalid_rom[  728] = 0; 
    i_addr_rom[  729] = 'h000006a0; 	    d_addr_rom[  729] = 'h00000f74; 	    wdata_rom[  729] = 'h9d5abb3e; 	    wvalid_rom[  729] = 0; 
    i_addr_rom[  730] = 'h00000290; 	    d_addr_rom[  730] = 'h00000fc0; 	    wdata_rom[  730] = 'hd74da7b2; 	    wvalid_rom[  730] = 0; 
    i_addr_rom[  731] = 'h00000404; 	    d_addr_rom[  731] = 'h00000c64; 	    wdata_rom[  731] = 'h8f152570; 	    wvalid_rom[  731] = 1; 
    i_addr_rom[  732] = 'h0000044c; 	    d_addr_rom[  732] = 'h00000d1c; 	    wdata_rom[  732] = 'h4cfe90e0; 	    wvalid_rom[  732] = 1; 
    i_addr_rom[  733] = 'h00000000; 	    d_addr_rom[  733] = 'h00000e60; 	    wdata_rom[  733] = 'h3434b45c; 	    wvalid_rom[  733] = 0; 
    i_addr_rom[  734] = 'h000000e8; 	    d_addr_rom[  734] = 'h00000f3c; 	    wdata_rom[  734] = 'h324f1e88; 	    wvalid_rom[  734] = 0; 
    i_addr_rom[  735] = 'h000003fc; 	    d_addr_rom[  735] = 'h00000fdc; 	    wdata_rom[  735] = 'h48be7dbc; 	    wvalid_rom[  735] = 0; 
    i_addr_rom[  736] = 'h00000330; 	    d_addr_rom[  736] = 'h00000a88; 	    wdata_rom[  736] = 'hd62e072f; 	    wvalid_rom[  736] = 1; 
    i_addr_rom[  737] = 'h00000228; 	    d_addr_rom[  737] = 'h00000b8c; 	    wdata_rom[  737] = 'h508d687c; 	    wvalid_rom[  737] = 0; 
    i_addr_rom[  738] = 'h000005e0; 	    d_addr_rom[  738] = 'h00000d38; 	    wdata_rom[  738] = 'hfd10760d; 	    wvalid_rom[  738] = 0; 
    i_addr_rom[  739] = 'h000001ec; 	    d_addr_rom[  739] = 'h00000e4c; 	    wdata_rom[  739] = 'h6c2c0112; 	    wvalid_rom[  739] = 1; 
    i_addr_rom[  740] = 'h00000068; 	    d_addr_rom[  740] = 'h00000b2c; 	    wdata_rom[  740] = 'h98dbd53e; 	    wvalid_rom[  740] = 1; 
    i_addr_rom[  741] = 'h00000648; 	    d_addr_rom[  741] = 'h00000b60; 	    wdata_rom[  741] = 'hd633445d; 	    wvalid_rom[  741] = 1; 
    i_addr_rom[  742] = 'h000000ac; 	    d_addr_rom[  742] = 'h00000e14; 	    wdata_rom[  742] = 'hb197c4a4; 	    wvalid_rom[  742] = 0; 
    i_addr_rom[  743] = 'h00000220; 	    d_addr_rom[  743] = 'h0000086c; 	    wdata_rom[  743] = 'h06b8a61e; 	    wvalid_rom[  743] = 0; 
    i_addr_rom[  744] = 'h00000560; 	    d_addr_rom[  744] = 'h00000934; 	    wdata_rom[  744] = 'h6a41a90d; 	    wvalid_rom[  744] = 0; 
    i_addr_rom[  745] = 'h00000394; 	    d_addr_rom[  745] = 'h00000c24; 	    wdata_rom[  745] = 'h4685f9a4; 	    wvalid_rom[  745] = 0; 
    i_addr_rom[  746] = 'h00000364; 	    d_addr_rom[  746] = 'h00000e20; 	    wdata_rom[  746] = 'ha417df24; 	    wvalid_rom[  746] = 1; 
    i_addr_rom[  747] = 'h000007f8; 	    d_addr_rom[  747] = 'h00000d98; 	    wdata_rom[  747] = 'hc480fc65; 	    wvalid_rom[  747] = 1; 
    i_addr_rom[  748] = 'h00000360; 	    d_addr_rom[  748] = 'h00000a40; 	    wdata_rom[  748] = 'hdbf35e38; 	    wvalid_rom[  748] = 0; 
    i_addr_rom[  749] = 'h00000338; 	    d_addr_rom[  749] = 'h00000c18; 	    wdata_rom[  749] = 'hbe05f5b5; 	    wvalid_rom[  749] = 1; 
    i_addr_rom[  750] = 'h00000668; 	    d_addr_rom[  750] = 'h00000db8; 	    wdata_rom[  750] = 'h0cefaeff; 	    wvalid_rom[  750] = 0; 
    i_addr_rom[  751] = 'h0000058c; 	    d_addr_rom[  751] = 'h00000a64; 	    wdata_rom[  751] = 'hf2fd5791; 	    wvalid_rom[  751] = 0; 
    i_addr_rom[  752] = 'h000004a8; 	    d_addr_rom[  752] = 'h000008d0; 	    wdata_rom[  752] = 'h549eecd2; 	    wvalid_rom[  752] = 0; 
    i_addr_rom[  753] = 'h000005ec; 	    d_addr_rom[  753] = 'h00000a30; 	    wdata_rom[  753] = 'hc052dabb; 	    wvalid_rom[  753] = 1; 
    i_addr_rom[  754] = 'h00000134; 	    d_addr_rom[  754] = 'h00000e08; 	    wdata_rom[  754] = 'hc10b4701; 	    wvalid_rom[  754] = 1; 
    i_addr_rom[  755] = 'h000001c4; 	    d_addr_rom[  755] = 'h00000ab4; 	    wdata_rom[  755] = 'hb693f1a1; 	    wvalid_rom[  755] = 1; 
    i_addr_rom[  756] = 'h000003b0; 	    d_addr_rom[  756] = 'h00000f7c; 	    wdata_rom[  756] = 'h858ad6e3; 	    wvalid_rom[  756] = 0; 
    i_addr_rom[  757] = 'h00000740; 	    d_addr_rom[  757] = 'h00000dac; 	    wdata_rom[  757] = 'hdd27f92d; 	    wvalid_rom[  757] = 1; 
    i_addr_rom[  758] = 'h000007f8; 	    d_addr_rom[  758] = 'h000009bc; 	    wdata_rom[  758] = 'h1d08eced; 	    wvalid_rom[  758] = 1; 
    i_addr_rom[  759] = 'h00000268; 	    d_addr_rom[  759] = 'h0000094c; 	    wdata_rom[  759] = 'hc6a133dd; 	    wvalid_rom[  759] = 1; 
    i_addr_rom[  760] = 'h0000066c; 	    d_addr_rom[  760] = 'h00000c4c; 	    wdata_rom[  760] = 'he4f21860; 	    wvalid_rom[  760] = 0; 
    i_addr_rom[  761] = 'h00000078; 	    d_addr_rom[  761] = 'h00000ef4; 	    wdata_rom[  761] = 'hca2940ec; 	    wvalid_rom[  761] = 0; 
    i_addr_rom[  762] = 'h00000170; 	    d_addr_rom[  762] = 'h00000bd0; 	    wdata_rom[  762] = 'h59e35b40; 	    wvalid_rom[  762] = 1; 
    i_addr_rom[  763] = 'h000001b4; 	    d_addr_rom[  763] = 'h00000bc8; 	    wdata_rom[  763] = 'h7c440eb8; 	    wvalid_rom[  763] = 0; 
    i_addr_rom[  764] = 'h00000414; 	    d_addr_rom[  764] = 'h00000cac; 	    wdata_rom[  764] = 'h7bea1e88; 	    wvalid_rom[  764] = 1; 
    i_addr_rom[  765] = 'h000002ac; 	    d_addr_rom[  765] = 'h000008f4; 	    wdata_rom[  765] = 'hfd137bc2; 	    wvalid_rom[  765] = 1; 
    i_addr_rom[  766] = 'h000002e8; 	    d_addr_rom[  766] = 'h00000904; 	    wdata_rom[  766] = 'h92a23d0f; 	    wvalid_rom[  766] = 0; 
    i_addr_rom[  767] = 'h00000644; 	    d_addr_rom[  767] = 'h00000cac; 	    wdata_rom[  767] = 'h2886db62; 	    wvalid_rom[  767] = 1; 
    i_addr_rom[  768] = 'h00000388; 	    d_addr_rom[  768] = 'h00000b98; 	    wdata_rom[  768] = 'hfb89ae4b; 	    wvalid_rom[  768] = 0; 
    i_addr_rom[  769] = 'h000000a4; 	    d_addr_rom[  769] = 'h00000a8c; 	    wdata_rom[  769] = 'hfa3e7336; 	    wvalid_rom[  769] = 1; 
    i_addr_rom[  770] = 'h000006c4; 	    d_addr_rom[  770] = 'h000008b0; 	    wdata_rom[  770] = 'h2ad11a7c; 	    wvalid_rom[  770] = 1; 
    i_addr_rom[  771] = 'h000001cc; 	    d_addr_rom[  771] = 'h00000d58; 	    wdata_rom[  771] = 'h43bfea76; 	    wvalid_rom[  771] = 1; 
    i_addr_rom[  772] = 'h00000364; 	    d_addr_rom[  772] = 'h00000dd4; 	    wdata_rom[  772] = 'h3c0ff2bc; 	    wvalid_rom[  772] = 0; 
    i_addr_rom[  773] = 'h00000168; 	    d_addr_rom[  773] = 'h00000d38; 	    wdata_rom[  773] = 'h7d778bf5; 	    wvalid_rom[  773] = 0; 
    i_addr_rom[  774] = 'h00000644; 	    d_addr_rom[  774] = 'h00000828; 	    wdata_rom[  774] = 'h3c85df91; 	    wvalid_rom[  774] = 1; 
    i_addr_rom[  775] = 'h00000704; 	    d_addr_rom[  775] = 'h00000d20; 	    wdata_rom[  775] = 'h1f88094c; 	    wvalid_rom[  775] = 0; 
    i_addr_rom[  776] = 'h000001ac; 	    d_addr_rom[  776] = 'h000008ec; 	    wdata_rom[  776] = 'h47b6a1d0; 	    wvalid_rom[  776] = 0; 
    i_addr_rom[  777] = 'h000002e0; 	    d_addr_rom[  777] = 'h00000a8c; 	    wdata_rom[  777] = 'h256d63e1; 	    wvalid_rom[  777] = 0; 
    i_addr_rom[  778] = 'h00000498; 	    d_addr_rom[  778] = 'h00000f30; 	    wdata_rom[  778] = 'h0f084ab1; 	    wvalid_rom[  778] = 1; 
    i_addr_rom[  779] = 'h000005ec; 	    d_addr_rom[  779] = 'h00000838; 	    wdata_rom[  779] = 'h3f685f74; 	    wvalid_rom[  779] = 0; 
    i_addr_rom[  780] = 'h0000064c; 	    d_addr_rom[  780] = 'h00000b04; 	    wdata_rom[  780] = 'h6c74bf7f; 	    wvalid_rom[  780] = 0; 
    i_addr_rom[  781] = 'h00000058; 	    d_addr_rom[  781] = 'h00000eb0; 	    wdata_rom[  781] = 'h72bb6c27; 	    wvalid_rom[  781] = 0; 
    i_addr_rom[  782] = 'h0000077c; 	    d_addr_rom[  782] = 'h00000d58; 	    wdata_rom[  782] = 'h7ba31f99; 	    wvalid_rom[  782] = 0; 
    i_addr_rom[  783] = 'h000000bc; 	    d_addr_rom[  783] = 'h00000b78; 	    wdata_rom[  783] = 'h1118f053; 	    wvalid_rom[  783] = 0; 
    i_addr_rom[  784] = 'h0000045c; 	    d_addr_rom[  784] = 'h00000908; 	    wdata_rom[  784] = 'h7a7ba5e4; 	    wvalid_rom[  784] = 0; 
    i_addr_rom[  785] = 'h000003ac; 	    d_addr_rom[  785] = 'h000009e4; 	    wdata_rom[  785] = 'h41519291; 	    wvalid_rom[  785] = 0; 
    i_addr_rom[  786] = 'h000006fc; 	    d_addr_rom[  786] = 'h00000b40; 	    wdata_rom[  786] = 'h63780c73; 	    wvalid_rom[  786] = 1; 
    i_addr_rom[  787] = 'h000007e4; 	    d_addr_rom[  787] = 'h00000aec; 	    wdata_rom[  787] = 'hdb76b6c5; 	    wvalid_rom[  787] = 0; 
    i_addr_rom[  788] = 'h000005c8; 	    d_addr_rom[  788] = 'h00000c24; 	    wdata_rom[  788] = 'h152a7194; 	    wvalid_rom[  788] = 0; 
    i_addr_rom[  789] = 'h00000634; 	    d_addr_rom[  789] = 'h00000a28; 	    wdata_rom[  789] = 'h5c5988ad; 	    wvalid_rom[  789] = 0; 
    i_addr_rom[  790] = 'h00000760; 	    d_addr_rom[  790] = 'h00000e7c; 	    wdata_rom[  790] = 'hae7148f9; 	    wvalid_rom[  790] = 0; 
    i_addr_rom[  791] = 'h000001fc; 	    d_addr_rom[  791] = 'h00000e4c; 	    wdata_rom[  791] = 'hc38ea955; 	    wvalid_rom[  791] = 1; 
    i_addr_rom[  792] = 'h00000158; 	    d_addr_rom[  792] = 'h00000b8c; 	    wdata_rom[  792] = 'hfe946c2c; 	    wvalid_rom[  792] = 1; 
    i_addr_rom[  793] = 'h0000066c; 	    d_addr_rom[  793] = 'h00000e98; 	    wdata_rom[  793] = 'h2dd82932; 	    wvalid_rom[  793] = 0; 
    i_addr_rom[  794] = 'h000005b0; 	    d_addr_rom[  794] = 'h000009d0; 	    wdata_rom[  794] = 'hea8fe672; 	    wvalid_rom[  794] = 1; 
    i_addr_rom[  795] = 'h000000d4; 	    d_addr_rom[  795] = 'h00000ae8; 	    wdata_rom[  795] = 'hbe04e2fe; 	    wvalid_rom[  795] = 0; 
    i_addr_rom[  796] = 'h000007f0; 	    d_addr_rom[  796] = 'h00000fe4; 	    wdata_rom[  796] = 'h031dac9d; 	    wvalid_rom[  796] = 1; 
    i_addr_rom[  797] = 'h00000568; 	    d_addr_rom[  797] = 'h00000ef4; 	    wdata_rom[  797] = 'hcc6d3967; 	    wvalid_rom[  797] = 1; 
    i_addr_rom[  798] = 'h0000031c; 	    d_addr_rom[  798] = 'h00000e80; 	    wdata_rom[  798] = 'h89d1289e; 	    wvalid_rom[  798] = 0; 
    i_addr_rom[  799] = 'h000000d0; 	    d_addr_rom[  799] = 'h00000bfc; 	    wdata_rom[  799] = 'h31fe316b; 	    wvalid_rom[  799] = 0; 
    i_addr_rom[  800] = 'h00000138; 	    d_addr_rom[  800] = 'h00000b50; 	    wdata_rom[  800] = 'hdb28f4b9; 	    wvalid_rom[  800] = 0; 
    i_addr_rom[  801] = 'h00000600; 	    d_addr_rom[  801] = 'h00000ef0; 	    wdata_rom[  801] = 'h617caffc; 	    wvalid_rom[  801] = 1; 
    i_addr_rom[  802] = 'h0000052c; 	    d_addr_rom[  802] = 'h00000bac; 	    wdata_rom[  802] = 'hc6df05c7; 	    wvalid_rom[  802] = 0; 
    i_addr_rom[  803] = 'h00000504; 	    d_addr_rom[  803] = 'h00000bb4; 	    wdata_rom[  803] = 'hbe084420; 	    wvalid_rom[  803] = 1; 
    i_addr_rom[  804] = 'h000004f8; 	    d_addr_rom[  804] = 'h000009bc; 	    wdata_rom[  804] = 'h8cf79887; 	    wvalid_rom[  804] = 1; 
    i_addr_rom[  805] = 'h000004bc; 	    d_addr_rom[  805] = 'h00000d4c; 	    wdata_rom[  805] = 'hca651fa1; 	    wvalid_rom[  805] = 0; 
    i_addr_rom[  806] = 'h000004dc; 	    d_addr_rom[  806] = 'h00000f64; 	    wdata_rom[  806] = 'ha0deaa6e; 	    wvalid_rom[  806] = 1; 
    i_addr_rom[  807] = 'h000004c8; 	    d_addr_rom[  807] = 'h0000083c; 	    wdata_rom[  807] = 'hdbef02e3; 	    wvalid_rom[  807] = 0; 
    i_addr_rom[  808] = 'h00000598; 	    d_addr_rom[  808] = 'h00000dcc; 	    wdata_rom[  808] = 'hb23e4793; 	    wvalid_rom[  808] = 1; 
    i_addr_rom[  809] = 'h000006f0; 	    d_addr_rom[  809] = 'h00000f98; 	    wdata_rom[  809] = 'h6f86f116; 	    wvalid_rom[  809] = 0; 
    i_addr_rom[  810] = 'h000003bc; 	    d_addr_rom[  810] = 'h00000b18; 	    wdata_rom[  810] = 'he94586c4; 	    wvalid_rom[  810] = 0; 
    i_addr_rom[  811] = 'h000000f0; 	    d_addr_rom[  811] = 'h00000910; 	    wdata_rom[  811] = 'h6fadf343; 	    wvalid_rom[  811] = 1; 
    i_addr_rom[  812] = 'h00000620; 	    d_addr_rom[  812] = 'h00000b40; 	    wdata_rom[  812] = 'h092da2a0; 	    wvalid_rom[  812] = 0; 
    i_addr_rom[  813] = 'h000001a0; 	    d_addr_rom[  813] = 'h000008e8; 	    wdata_rom[  813] = 'h3fd6ce0f; 	    wvalid_rom[  813] = 0; 
    i_addr_rom[  814] = 'h000000e0; 	    d_addr_rom[  814] = 'h00000fcc; 	    wdata_rom[  814] = 'h1e81152b; 	    wvalid_rom[  814] = 0; 
    i_addr_rom[  815] = 'h000006cc; 	    d_addr_rom[  815] = 'h000008dc; 	    wdata_rom[  815] = 'h88d95f23; 	    wvalid_rom[  815] = 1; 
    i_addr_rom[  816] = 'h00000050; 	    d_addr_rom[  816] = 'h00000f90; 	    wdata_rom[  816] = 'hc160ddfb; 	    wvalid_rom[  816] = 0; 
    i_addr_rom[  817] = 'h00000208; 	    d_addr_rom[  817] = 'h00000a00; 	    wdata_rom[  817] = 'h5c8e7e38; 	    wvalid_rom[  817] = 0; 
    i_addr_rom[  818] = 'h000007a8; 	    d_addr_rom[  818] = 'h00000f14; 	    wdata_rom[  818] = 'hb2ed62bb; 	    wvalid_rom[  818] = 1; 
    i_addr_rom[  819] = 'h000006b4; 	    d_addr_rom[  819] = 'h00000800; 	    wdata_rom[  819] = 'hf0ac6b0d; 	    wvalid_rom[  819] = 0; 
    i_addr_rom[  820] = 'h0000016c; 	    d_addr_rom[  820] = 'h00000d50; 	    wdata_rom[  820] = 'h171c925c; 	    wvalid_rom[  820] = 0; 
    i_addr_rom[  821] = 'h000000cc; 	    d_addr_rom[  821] = 'h00000c50; 	    wdata_rom[  821] = 'h4138d38f; 	    wvalid_rom[  821] = 1; 
    i_addr_rom[  822] = 'h000005a4; 	    d_addr_rom[  822] = 'h00000b54; 	    wdata_rom[  822] = 'h7735f1d7; 	    wvalid_rom[  822] = 1; 
    i_addr_rom[  823] = 'h0000046c; 	    d_addr_rom[  823] = 'h00000b2c; 	    wdata_rom[  823] = 'hcb17ed59; 	    wvalid_rom[  823] = 1; 
    i_addr_rom[  824] = 'h00000614; 	    d_addr_rom[  824] = 'h00000ca4; 	    wdata_rom[  824] = 'h776b66f4; 	    wvalid_rom[  824] = 0; 
    i_addr_rom[  825] = 'h000002ec; 	    d_addr_rom[  825] = 'h00000838; 	    wdata_rom[  825] = 'h1825a790; 	    wvalid_rom[  825] = 0; 
    i_addr_rom[  826] = 'h000006b4; 	    d_addr_rom[  826] = 'h00000a24; 	    wdata_rom[  826] = 'h2097e19b; 	    wvalid_rom[  826] = 1; 
    i_addr_rom[  827] = 'h00000060; 	    d_addr_rom[  827] = 'h00000c0c; 	    wdata_rom[  827] = 'hffa99abb; 	    wvalid_rom[  827] = 0; 
    i_addr_rom[  828] = 'h000005c0; 	    d_addr_rom[  828] = 'h00000e00; 	    wdata_rom[  828] = 'h798ef231; 	    wvalid_rom[  828] = 0; 
    i_addr_rom[  829] = 'h000002f4; 	    d_addr_rom[  829] = 'h00000e08; 	    wdata_rom[  829] = 'h2da1d663; 	    wvalid_rom[  829] = 1; 
    i_addr_rom[  830] = 'h000007f4; 	    d_addr_rom[  830] = 'h00000cb4; 	    wdata_rom[  830] = 'h48e69460; 	    wvalid_rom[  830] = 0; 
    i_addr_rom[  831] = 'h000006f4; 	    d_addr_rom[  831] = 'h00000cf0; 	    wdata_rom[  831] = 'ha78c6993; 	    wvalid_rom[  831] = 0; 
    i_addr_rom[  832] = 'h00000348; 	    d_addr_rom[  832] = 'h00000e64; 	    wdata_rom[  832] = 'hf6573af3; 	    wvalid_rom[  832] = 0; 
    i_addr_rom[  833] = 'h0000020c; 	    d_addr_rom[  833] = 'h00000e00; 	    wdata_rom[  833] = 'h5b1335f3; 	    wvalid_rom[  833] = 1; 
    i_addr_rom[  834] = 'h000006f0; 	    d_addr_rom[  834] = 'h00000a68; 	    wdata_rom[  834] = 'h7b83487f; 	    wvalid_rom[  834] = 1; 
    i_addr_rom[  835] = 'h00000074; 	    d_addr_rom[  835] = 'h00000f0c; 	    wdata_rom[  835] = 'hf99d6ed4; 	    wvalid_rom[  835] = 1; 
    i_addr_rom[  836] = 'h00000178; 	    d_addr_rom[  836] = 'h00000b38; 	    wdata_rom[  836] = 'h11d67291; 	    wvalid_rom[  836] = 1; 
    i_addr_rom[  837] = 'h000001cc; 	    d_addr_rom[  837] = 'h00000bdc; 	    wdata_rom[  837] = 'h1b34be14; 	    wvalid_rom[  837] = 0; 
    i_addr_rom[  838] = 'h000002dc; 	    d_addr_rom[  838] = 'h00000a88; 	    wdata_rom[  838] = 'h3cfebba7; 	    wvalid_rom[  838] = 1; 
    i_addr_rom[  839] = 'h0000013c; 	    d_addr_rom[  839] = 'h00000934; 	    wdata_rom[  839] = 'hf4991051; 	    wvalid_rom[  839] = 1; 
    i_addr_rom[  840] = 'h00000420; 	    d_addr_rom[  840] = 'h00000f48; 	    wdata_rom[  840] = 'h9872f292; 	    wvalid_rom[  840] = 1; 
    i_addr_rom[  841] = 'h000007f8; 	    d_addr_rom[  841] = 'h00000c38; 	    wdata_rom[  841] = 'h2de8ec03; 	    wvalid_rom[  841] = 1; 
    i_addr_rom[  842] = 'h0000020c; 	    d_addr_rom[  842] = 'h00000a80; 	    wdata_rom[  842] = 'hfa4fb743; 	    wvalid_rom[  842] = 0; 
    i_addr_rom[  843] = 'h00000184; 	    d_addr_rom[  843] = 'h00000cb4; 	    wdata_rom[  843] = 'h373a9814; 	    wvalid_rom[  843] = 1; 
    i_addr_rom[  844] = 'h000002d0; 	    d_addr_rom[  844] = 'h00000e08; 	    wdata_rom[  844] = 'h8a1cd289; 	    wvalid_rom[  844] = 0; 
    i_addr_rom[  845] = 'h00000314; 	    d_addr_rom[  845] = 'h00000aa8; 	    wdata_rom[  845] = 'h64934c12; 	    wvalid_rom[  845] = 1; 
    i_addr_rom[  846] = 'h000000cc; 	    d_addr_rom[  846] = 'h00000f38; 	    wdata_rom[  846] = 'h5a10d2ea; 	    wvalid_rom[  846] = 0; 
    i_addr_rom[  847] = 'h00000774; 	    d_addr_rom[  847] = 'h000009e8; 	    wdata_rom[  847] = 'h575109f9; 	    wvalid_rom[  847] = 0; 
    i_addr_rom[  848] = 'h00000530; 	    d_addr_rom[  848] = 'h000009a8; 	    wdata_rom[  848] = 'h6bb34993; 	    wvalid_rom[  848] = 1; 
    i_addr_rom[  849] = 'h00000024; 	    d_addr_rom[  849] = 'h00000fa8; 	    wdata_rom[  849] = 'h492a9ea4; 	    wvalid_rom[  849] = 0; 
    i_addr_rom[  850] = 'h000005f4; 	    d_addr_rom[  850] = 'h00000c38; 	    wdata_rom[  850] = 'hb9e8a2c5; 	    wvalid_rom[  850] = 0; 
    i_addr_rom[  851] = 'h000007e8; 	    d_addr_rom[  851] = 'h00000d64; 	    wdata_rom[  851] = 'h42da9996; 	    wvalid_rom[  851] = 1; 
    i_addr_rom[  852] = 'h000005e0; 	    d_addr_rom[  852] = 'h00000ff4; 	    wdata_rom[  852] = 'h47d5a114; 	    wvalid_rom[  852] = 0; 
    i_addr_rom[  853] = 'h00000100; 	    d_addr_rom[  853] = 'h00000cb8; 	    wdata_rom[  853] = 'hde03ba82; 	    wvalid_rom[  853] = 0; 
    i_addr_rom[  854] = 'h000007e4; 	    d_addr_rom[  854] = 'h00000b2c; 	    wdata_rom[  854] = 'h1ce8d6fd; 	    wvalid_rom[  854] = 0; 
    i_addr_rom[  855] = 'h00000528; 	    d_addr_rom[  855] = 'h00000e48; 	    wdata_rom[  855] = 'h561aeda5; 	    wvalid_rom[  855] = 0; 
    i_addr_rom[  856] = 'h000006c4; 	    d_addr_rom[  856] = 'h00000f48; 	    wdata_rom[  856] = 'hc81d62e7; 	    wvalid_rom[  856] = 0; 
    i_addr_rom[  857] = 'h000006a8; 	    d_addr_rom[  857] = 'h000008b4; 	    wdata_rom[  857] = 'hfb6d07f4; 	    wvalid_rom[  857] = 1; 
    i_addr_rom[  858] = 'h00000788; 	    d_addr_rom[  858] = 'h00000878; 	    wdata_rom[  858] = 'h4e14e39c; 	    wvalid_rom[  858] = 0; 
    i_addr_rom[  859] = 'h000006b0; 	    d_addr_rom[  859] = 'h00000abc; 	    wdata_rom[  859] = 'hf300425e; 	    wvalid_rom[  859] = 1; 
    i_addr_rom[  860] = 'h000001a4; 	    d_addr_rom[  860] = 'h00000ac8; 	    wdata_rom[  860] = 'h7cd9f6c5; 	    wvalid_rom[  860] = 1; 
    i_addr_rom[  861] = 'h00000314; 	    d_addr_rom[  861] = 'h00000d90; 	    wdata_rom[  861] = 'h90350731; 	    wvalid_rom[  861] = 1; 
    i_addr_rom[  862] = 'h00000784; 	    d_addr_rom[  862] = 'h00000950; 	    wdata_rom[  862] = 'hecb20f8b; 	    wvalid_rom[  862] = 0; 
    i_addr_rom[  863] = 'h00000124; 	    d_addr_rom[  863] = 'h00000928; 	    wdata_rom[  863] = 'h6f9286ac; 	    wvalid_rom[  863] = 1; 
    i_addr_rom[  864] = 'h00000338; 	    d_addr_rom[  864] = 'h00000e90; 	    wdata_rom[  864] = 'hf6b684ad; 	    wvalid_rom[  864] = 0; 
    i_addr_rom[  865] = 'h00000288; 	    d_addr_rom[  865] = 'h00000978; 	    wdata_rom[  865] = 'h03aa106e; 	    wvalid_rom[  865] = 0; 
    i_addr_rom[  866] = 'h00000600; 	    d_addr_rom[  866] = 'h00000f90; 	    wdata_rom[  866] = 'h5179fb17; 	    wvalid_rom[  866] = 0; 
    i_addr_rom[  867] = 'h000007bc; 	    d_addr_rom[  867] = 'h00000f0c; 	    wdata_rom[  867] = 'hb816c594; 	    wvalid_rom[  867] = 0; 
    i_addr_rom[  868] = 'h00000430; 	    d_addr_rom[  868] = 'h00000ad8; 	    wdata_rom[  868] = 'h755c8395; 	    wvalid_rom[  868] = 1; 
    i_addr_rom[  869] = 'h000005d0; 	    d_addr_rom[  869] = 'h00000a04; 	    wdata_rom[  869] = 'hc673af60; 	    wvalid_rom[  869] = 0; 
    i_addr_rom[  870] = 'h000005c8; 	    d_addr_rom[  870] = 'h00000b8c; 	    wdata_rom[  870] = 'h3f48c082; 	    wvalid_rom[  870] = 0; 
    i_addr_rom[  871] = 'h00000158; 	    d_addr_rom[  871] = 'h00000b54; 	    wdata_rom[  871] = 'h5a1e46b9; 	    wvalid_rom[  871] = 0; 
    i_addr_rom[  872] = 'h00000160; 	    d_addr_rom[  872] = 'h000009cc; 	    wdata_rom[  872] = 'h688b8ebe; 	    wvalid_rom[  872] = 1; 
    i_addr_rom[  873] = 'h00000438; 	    d_addr_rom[  873] = 'h00000bdc; 	    wdata_rom[  873] = 'h57c4c1c4; 	    wvalid_rom[  873] = 1; 
    i_addr_rom[  874] = 'h000005a4; 	    d_addr_rom[  874] = 'h0000088c; 	    wdata_rom[  874] = 'hd99ee10e; 	    wvalid_rom[  874] = 1; 
    i_addr_rom[  875] = 'h00000350; 	    d_addr_rom[  875] = 'h00000de8; 	    wdata_rom[  875] = 'he4b7b24a; 	    wvalid_rom[  875] = 0; 
    i_addr_rom[  876] = 'h00000474; 	    d_addr_rom[  876] = 'h00000e74; 	    wdata_rom[  876] = 'h8d8e612f; 	    wvalid_rom[  876] = 1; 
    i_addr_rom[  877] = 'h000003e4; 	    d_addr_rom[  877] = 'h00000b50; 	    wdata_rom[  877] = 'hd17afea4; 	    wvalid_rom[  877] = 0; 
    i_addr_rom[  878] = 'h00000374; 	    d_addr_rom[  878] = 'h00000f84; 	    wdata_rom[  878] = 'hc0bc6993; 	    wvalid_rom[  878] = 1; 
    i_addr_rom[  879] = 'h00000094; 	    d_addr_rom[  879] = 'h00000be4; 	    wdata_rom[  879] = 'h8d218809; 	    wvalid_rom[  879] = 1; 
    i_addr_rom[  880] = 'h0000037c; 	    d_addr_rom[  880] = 'h00000ec0; 	    wdata_rom[  880] = 'h18b0bb8d; 	    wvalid_rom[  880] = 1; 
    i_addr_rom[  881] = 'h00000530; 	    d_addr_rom[  881] = 'h00000fdc; 	    wdata_rom[  881] = 'h8172b2ba; 	    wvalid_rom[  881] = 1; 
    i_addr_rom[  882] = 'h000004a8; 	    d_addr_rom[  882] = 'h0000086c; 	    wdata_rom[  882] = 'hc85c8e85; 	    wvalid_rom[  882] = 0; 
    i_addr_rom[  883] = 'h00000138; 	    d_addr_rom[  883] = 'h00000dd0; 	    wdata_rom[  883] = 'he4e7cdda; 	    wvalid_rom[  883] = 1; 
    i_addr_rom[  884] = 'h00000668; 	    d_addr_rom[  884] = 'h00000cbc; 	    wdata_rom[  884] = 'h3965efd2; 	    wvalid_rom[  884] = 0; 
    i_addr_rom[  885] = 'h000007c0; 	    d_addr_rom[  885] = 'h00000ee8; 	    wdata_rom[  885] = 'he0876766; 	    wvalid_rom[  885] = 0; 
    i_addr_rom[  886] = 'h000007e4; 	    d_addr_rom[  886] = 'h0000080c; 	    wdata_rom[  886] = 'h30ceef7e; 	    wvalid_rom[  886] = 1; 
    i_addr_rom[  887] = 'h0000069c; 	    d_addr_rom[  887] = 'h00000860; 	    wdata_rom[  887] = 'h07fd82c0; 	    wvalid_rom[  887] = 1; 
    i_addr_rom[  888] = 'h00000258; 	    d_addr_rom[  888] = 'h00000bfc; 	    wdata_rom[  888] = 'h8699c912; 	    wvalid_rom[  888] = 1; 
    i_addr_rom[  889] = 'h00000770; 	    d_addr_rom[  889] = 'h00000fa0; 	    wdata_rom[  889] = 'h10198418; 	    wvalid_rom[  889] = 1; 
    i_addr_rom[  890] = 'h00000078; 	    d_addr_rom[  890] = 'h00000d7c; 	    wdata_rom[  890] = 'hcc7b6666; 	    wvalid_rom[  890] = 1; 
    i_addr_rom[  891] = 'h000002a4; 	    d_addr_rom[  891] = 'h00000b24; 	    wdata_rom[  891] = 'hbe5ca57f; 	    wvalid_rom[  891] = 0; 
    i_addr_rom[  892] = 'h00000170; 	    d_addr_rom[  892] = 'h00000bf0; 	    wdata_rom[  892] = 'h03b149e1; 	    wvalid_rom[  892] = 0; 
    i_addr_rom[  893] = 'h00000104; 	    d_addr_rom[  893] = 'h00000c34; 	    wdata_rom[  893] = 'h62f0ed9e; 	    wvalid_rom[  893] = 0; 
    i_addr_rom[  894] = 'h000001c0; 	    d_addr_rom[  894] = 'h00000c74; 	    wdata_rom[  894] = 'hd7456174; 	    wvalid_rom[  894] = 0; 
    i_addr_rom[  895] = 'h00000154; 	    d_addr_rom[  895] = 'h00000cbc; 	    wdata_rom[  895] = 'h86a1b8f6; 	    wvalid_rom[  895] = 0; 
    i_addr_rom[  896] = 'h00000490; 	    d_addr_rom[  896] = 'h00000ed4; 	    wdata_rom[  896] = 'h5f529b49; 	    wvalid_rom[  896] = 0; 
    i_addr_rom[  897] = 'h00000714; 	    d_addr_rom[  897] = 'h00000a44; 	    wdata_rom[  897] = 'h25e20b2a; 	    wvalid_rom[  897] = 1; 
    i_addr_rom[  898] = 'h000002ec; 	    d_addr_rom[  898] = 'h00000e1c; 	    wdata_rom[  898] = 'hdd01bd8e; 	    wvalid_rom[  898] = 1; 
    i_addr_rom[  899] = 'h000000d0; 	    d_addr_rom[  899] = 'h00000a98; 	    wdata_rom[  899] = 'hc1e5200e; 	    wvalid_rom[  899] = 0; 
    i_addr_rom[  900] = 'h00000700; 	    d_addr_rom[  900] = 'h00000b48; 	    wdata_rom[  900] = 'h2514bee8; 	    wvalid_rom[  900] = 0; 
    i_addr_rom[  901] = 'h0000011c; 	    d_addr_rom[  901] = 'h00000b70; 	    wdata_rom[  901] = 'hd47aa980; 	    wvalid_rom[  901] = 0; 
    i_addr_rom[  902] = 'h00000274; 	    d_addr_rom[  902] = 'h00000904; 	    wdata_rom[  902] = 'he7891e0a; 	    wvalid_rom[  902] = 0; 
    i_addr_rom[  903] = 'h000005a8; 	    d_addr_rom[  903] = 'h00000ce8; 	    wdata_rom[  903] = 'hf89c7e83; 	    wvalid_rom[  903] = 0; 
    i_addr_rom[  904] = 'h000002c4; 	    d_addr_rom[  904] = 'h00000a58; 	    wdata_rom[  904] = 'h1cb7624b; 	    wvalid_rom[  904] = 0; 
    i_addr_rom[  905] = 'h0000059c; 	    d_addr_rom[  905] = 'h00000ed8; 	    wdata_rom[  905] = 'h54fa4c0e; 	    wvalid_rom[  905] = 1; 
    i_addr_rom[  906] = 'h0000051c; 	    d_addr_rom[  906] = 'h00000eac; 	    wdata_rom[  906] = 'hd8f175a3; 	    wvalid_rom[  906] = 0; 
    i_addr_rom[  907] = 'h000005b4; 	    d_addr_rom[  907] = 'h00000d78; 	    wdata_rom[  907] = 'h1d139616; 	    wvalid_rom[  907] = 1; 
    i_addr_rom[  908] = 'h000004e0; 	    d_addr_rom[  908] = 'h00000ddc; 	    wdata_rom[  908] = 'hfb9502ed; 	    wvalid_rom[  908] = 1; 
    i_addr_rom[  909] = 'h00000234; 	    d_addr_rom[  909] = 'h00000a44; 	    wdata_rom[  909] = 'hec519282; 	    wvalid_rom[  909] = 1; 
    i_addr_rom[  910] = 'h000005d4; 	    d_addr_rom[  910] = 'h00000d70; 	    wdata_rom[  910] = 'h38aa525f; 	    wvalid_rom[  910] = 1; 
    i_addr_rom[  911] = 'h000006c8; 	    d_addr_rom[  911] = 'h00000aa0; 	    wdata_rom[  911] = 'hf3800c81; 	    wvalid_rom[  911] = 0; 
    i_addr_rom[  912] = 'h000000d8; 	    d_addr_rom[  912] = 'h00000de4; 	    wdata_rom[  912] = 'h1fcb94fc; 	    wvalid_rom[  912] = 1; 
    i_addr_rom[  913] = 'h00000680; 	    d_addr_rom[  913] = 'h00000a3c; 	    wdata_rom[  913] = 'h4c14dcfd; 	    wvalid_rom[  913] = 0; 
    i_addr_rom[  914] = 'h00000130; 	    d_addr_rom[  914] = 'h0000094c; 	    wdata_rom[  914] = 'he10f5652; 	    wvalid_rom[  914] = 1; 
    i_addr_rom[  915] = 'h000001c0; 	    d_addr_rom[  915] = 'h00000e68; 	    wdata_rom[  915] = 'hf953444d; 	    wvalid_rom[  915] = 0; 
    i_addr_rom[  916] = 'h000000ac; 	    d_addr_rom[  916] = 'h00000abc; 	    wdata_rom[  916] = 'h3b3dbacf; 	    wvalid_rom[  916] = 0; 
    i_addr_rom[  917] = 'h000006a0; 	    d_addr_rom[  917] = 'h00000830; 	    wdata_rom[  917] = 'h3ce07fb1; 	    wvalid_rom[  917] = 0; 
    i_addr_rom[  918] = 'h00000538; 	    d_addr_rom[  918] = 'h000009c4; 	    wdata_rom[  918] = 'hc33ee94c; 	    wvalid_rom[  918] = 0; 
    i_addr_rom[  919] = 'h000006d8; 	    d_addr_rom[  919] = 'h00000a94; 	    wdata_rom[  919] = 'hcd03d0f0; 	    wvalid_rom[  919] = 0; 
    i_addr_rom[  920] = 'h00000414; 	    d_addr_rom[  920] = 'h00000cb0; 	    wdata_rom[  920] = 'h536382ac; 	    wvalid_rom[  920] = 0; 
    i_addr_rom[  921] = 'h00000304; 	    d_addr_rom[  921] = 'h00000980; 	    wdata_rom[  921] = 'h4d2114c3; 	    wvalid_rom[  921] = 0; 
    i_addr_rom[  922] = 'h000002d0; 	    d_addr_rom[  922] = 'h0000098c; 	    wdata_rom[  922] = 'hcb2dd2d5; 	    wvalid_rom[  922] = 1; 
    i_addr_rom[  923] = 'h00000200; 	    d_addr_rom[  923] = 'h00000cb8; 	    wdata_rom[  923] = 'h76e869dc; 	    wvalid_rom[  923] = 0; 
    i_addr_rom[  924] = 'h0000053c; 	    d_addr_rom[  924] = 'h00000d70; 	    wdata_rom[  924] = 'h0f0d3218; 	    wvalid_rom[  924] = 0; 
    i_addr_rom[  925] = 'h000001fc; 	    d_addr_rom[  925] = 'h00000c80; 	    wdata_rom[  925] = 'hbbe74d81; 	    wvalid_rom[  925] = 1; 
    i_addr_rom[  926] = 'h000000e0; 	    d_addr_rom[  926] = 'h00000ae8; 	    wdata_rom[  926] = 'h9f980a01; 	    wvalid_rom[  926] = 0; 
    i_addr_rom[  927] = 'h000002a8; 	    d_addr_rom[  927] = 'h00000d78; 	    wdata_rom[  927] = 'hc89a791f; 	    wvalid_rom[  927] = 1; 
    i_addr_rom[  928] = 'h000001d0; 	    d_addr_rom[  928] = 'h00000878; 	    wdata_rom[  928] = 'h5768c071; 	    wvalid_rom[  928] = 1; 
    i_addr_rom[  929] = 'h00000564; 	    d_addr_rom[  929] = 'h00000c78; 	    wdata_rom[  929] = 'h85709fbf; 	    wvalid_rom[  929] = 0; 
    i_addr_rom[  930] = 'h000005f4; 	    d_addr_rom[  930] = 'h00000ce4; 	    wdata_rom[  930] = 'h24512bcb; 	    wvalid_rom[  930] = 0; 
    i_addr_rom[  931] = 'h00000650; 	    d_addr_rom[  931] = 'h00000808; 	    wdata_rom[  931] = 'hd6220b67; 	    wvalid_rom[  931] = 0; 
    i_addr_rom[  932] = 'h000005d4; 	    d_addr_rom[  932] = 'h00000ed4; 	    wdata_rom[  932] = 'h471cb4db; 	    wvalid_rom[  932] = 1; 
    i_addr_rom[  933] = 'h00000154; 	    d_addr_rom[  933] = 'h00000a88; 	    wdata_rom[  933] = 'h8dbe5573; 	    wvalid_rom[  933] = 0; 
    i_addr_rom[  934] = 'h00000538; 	    d_addr_rom[  934] = 'h00000f18; 	    wdata_rom[  934] = 'h6fb136a9; 	    wvalid_rom[  934] = 1; 
    i_addr_rom[  935] = 'h00000474; 	    d_addr_rom[  935] = 'h00000e64; 	    wdata_rom[  935] = 'h8681b020; 	    wvalid_rom[  935] = 0; 
    i_addr_rom[  936] = 'h000002ac; 	    d_addr_rom[  936] = 'h000009ac; 	    wdata_rom[  936] = 'hdc0275fb; 	    wvalid_rom[  936] = 1; 
    i_addr_rom[  937] = 'h0000034c; 	    d_addr_rom[  937] = 'h00000f00; 	    wdata_rom[  937] = 'hee16184b; 	    wvalid_rom[  937] = 0; 
    i_addr_rom[  938] = 'h000004c4; 	    d_addr_rom[  938] = 'h00000cb0; 	    wdata_rom[  938] = 'hf7a76e2b; 	    wvalid_rom[  938] = 0; 
    i_addr_rom[  939] = 'h00000174; 	    d_addr_rom[  939] = 'h00000810; 	    wdata_rom[  939] = 'hbc4f5bfd; 	    wvalid_rom[  939] = 1; 
    i_addr_rom[  940] = 'h0000011c; 	    d_addr_rom[  940] = 'h00000bc8; 	    wdata_rom[  940] = 'h22b91f48; 	    wvalid_rom[  940] = 1; 
    i_addr_rom[  941] = 'h0000070c; 	    d_addr_rom[  941] = 'h00000b9c; 	    wdata_rom[  941] = 'h21634f23; 	    wvalid_rom[  941] = 1; 
    i_addr_rom[  942] = 'h00000500; 	    d_addr_rom[  942] = 'h0000088c; 	    wdata_rom[  942] = 'hf171825b; 	    wvalid_rom[  942] = 0; 
    i_addr_rom[  943] = 'h000000e8; 	    d_addr_rom[  943] = 'h00000ad8; 	    wdata_rom[  943] = 'hd08ee915; 	    wvalid_rom[  943] = 1; 
    i_addr_rom[  944] = 'h000006a4; 	    d_addr_rom[  944] = 'h00000e28; 	    wdata_rom[  944] = 'h597898d7; 	    wvalid_rom[  944] = 1; 
    i_addr_rom[  945] = 'h000003a4; 	    d_addr_rom[  945] = 'h0000085c; 	    wdata_rom[  945] = 'hfa4cd90f; 	    wvalid_rom[  945] = 0; 
    i_addr_rom[  946] = 'h000001ac; 	    d_addr_rom[  946] = 'h00000cf4; 	    wdata_rom[  946] = 'h09f1e248; 	    wvalid_rom[  946] = 1; 
    i_addr_rom[  947] = 'h00000704; 	    d_addr_rom[  947] = 'h00000968; 	    wdata_rom[  947] = 'h4e2ddc2b; 	    wvalid_rom[  947] = 1; 
    i_addr_rom[  948] = 'h000000c4; 	    d_addr_rom[  948] = 'h00000dc0; 	    wdata_rom[  948] = 'hfc36d05c; 	    wvalid_rom[  948] = 0; 
    i_addr_rom[  949] = 'h0000032c; 	    d_addr_rom[  949] = 'h00000f74; 	    wdata_rom[  949] = 'hba8fd2f6; 	    wvalid_rom[  949] = 0; 
    i_addr_rom[  950] = 'h000006cc; 	    d_addr_rom[  950] = 'h00000dd0; 	    wdata_rom[  950] = 'h3d9fc0ef; 	    wvalid_rom[  950] = 0; 
    i_addr_rom[  951] = 'h000007a8; 	    d_addr_rom[  951] = 'h00000fd8; 	    wdata_rom[  951] = 'h2040b654; 	    wvalid_rom[  951] = 1; 
    i_addr_rom[  952] = 'h00000414; 	    d_addr_rom[  952] = 'h00000f6c; 	    wdata_rom[  952] = 'hcb63c8fe; 	    wvalid_rom[  952] = 0; 
    i_addr_rom[  953] = 'h000000c0; 	    d_addr_rom[  953] = 'h0000087c; 	    wdata_rom[  953] = 'h6a21edef; 	    wvalid_rom[  953] = 1; 
    i_addr_rom[  954] = 'h000001bc; 	    d_addr_rom[  954] = 'h00000dec; 	    wdata_rom[  954] = 'h3c3b96d5; 	    wvalid_rom[  954] = 1; 
    i_addr_rom[  955] = 'h00000260; 	    d_addr_rom[  955] = 'h00000bac; 	    wdata_rom[  955] = 'h50459330; 	    wvalid_rom[  955] = 0; 
    i_addr_rom[  956] = 'h00000790; 	    d_addr_rom[  956] = 'h000008f8; 	    wdata_rom[  956] = 'hbfd1c8bd; 	    wvalid_rom[  956] = 0; 
    i_addr_rom[  957] = 'h000001d8; 	    d_addr_rom[  957] = 'h00000de8; 	    wdata_rom[  957] = 'ha8820b0a; 	    wvalid_rom[  957] = 0; 
    i_addr_rom[  958] = 'h00000394; 	    d_addr_rom[  958] = 'h00000e14; 	    wdata_rom[  958] = 'h4640ef05; 	    wvalid_rom[  958] = 0; 
    i_addr_rom[  959] = 'h0000006c; 	    d_addr_rom[  959] = 'h00000800; 	    wdata_rom[  959] = 'h2d1f69dc; 	    wvalid_rom[  959] = 0; 
    i_addr_rom[  960] = 'h00000584; 	    d_addr_rom[  960] = 'h00000e3c; 	    wdata_rom[  960] = 'h38af5f05; 	    wvalid_rom[  960] = 0; 
    i_addr_rom[  961] = 'h00000094; 	    d_addr_rom[  961] = 'h00000a98; 	    wdata_rom[  961] = 'h1f69f6cd; 	    wvalid_rom[  961] = 1; 
    i_addr_rom[  962] = 'h00000324; 	    d_addr_rom[  962] = 'h00000c2c; 	    wdata_rom[  962] = 'he8b0ca7f; 	    wvalid_rom[  962] = 0; 
    i_addr_rom[  963] = 'h000007a8; 	    d_addr_rom[  963] = 'h00000dd8; 	    wdata_rom[  963] = 'hf704bc80; 	    wvalid_rom[  963] = 0; 
    i_addr_rom[  964] = 'h000003dc; 	    d_addr_rom[  964] = 'h00000a68; 	    wdata_rom[  964] = 'hdab8d48e; 	    wvalid_rom[  964] = 0; 
    i_addr_rom[  965] = 'h00000528; 	    d_addr_rom[  965] = 'h00000844; 	    wdata_rom[  965] = 'h79420320; 	    wvalid_rom[  965] = 0; 
    i_addr_rom[  966] = 'h00000488; 	    d_addr_rom[  966] = 'h00000914; 	    wdata_rom[  966] = 'h0bdb6e26; 	    wvalid_rom[  966] = 0; 
    i_addr_rom[  967] = 'h00000274; 	    d_addr_rom[  967] = 'h00000a44; 	    wdata_rom[  967] = 'hfc2d4c34; 	    wvalid_rom[  967] = 0; 
    i_addr_rom[  968] = 'h00000614; 	    d_addr_rom[  968] = 'h000009d4; 	    wdata_rom[  968] = 'h9e478c3d; 	    wvalid_rom[  968] = 0; 
    i_addr_rom[  969] = 'h000005f0; 	    d_addr_rom[  969] = 'h00000d08; 	    wdata_rom[  969] = 'h0d0a0e11; 	    wvalid_rom[  969] = 0; 
    i_addr_rom[  970] = 'h000001bc; 	    d_addr_rom[  970] = 'h00000918; 	    wdata_rom[  970] = 'h87b8ca4b; 	    wvalid_rom[  970] = 1; 
    i_addr_rom[  971] = 'h00000484; 	    d_addr_rom[  971] = 'h00000e98; 	    wdata_rom[  971] = 'hd26b9b17; 	    wvalid_rom[  971] = 1; 
    i_addr_rom[  972] = 'h00000330; 	    d_addr_rom[  972] = 'h00000f98; 	    wdata_rom[  972] = 'h206119af; 	    wvalid_rom[  972] = 0; 
    i_addr_rom[  973] = 'h00000198; 	    d_addr_rom[  973] = 'h00000c64; 	    wdata_rom[  973] = 'ha40513b6; 	    wvalid_rom[  973] = 1; 
    i_addr_rom[  974] = 'h00000078; 	    d_addr_rom[  974] = 'h00000bd4; 	    wdata_rom[  974] = 'h4478bfc0; 	    wvalid_rom[  974] = 1; 
    i_addr_rom[  975] = 'h00000460; 	    d_addr_rom[  975] = 'h00000f18; 	    wdata_rom[  975] = 'h68f91cea; 	    wvalid_rom[  975] = 0; 
    i_addr_rom[  976] = 'h00000750; 	    d_addr_rom[  976] = 'h00000a44; 	    wdata_rom[  976] = 'hd66e2cc4; 	    wvalid_rom[  976] = 1; 
    i_addr_rom[  977] = 'h0000067c; 	    d_addr_rom[  977] = 'h00000f30; 	    wdata_rom[  977] = 'h5ef6c847; 	    wvalid_rom[  977] = 1; 
    i_addr_rom[  978] = 'h00000494; 	    d_addr_rom[  978] = 'h00000d10; 	    wdata_rom[  978] = 'h898b4ae9; 	    wvalid_rom[  978] = 1; 
    i_addr_rom[  979] = 'h00000280; 	    d_addr_rom[  979] = 'h000009b8; 	    wdata_rom[  979] = 'h3427832b; 	    wvalid_rom[  979] = 1; 
    i_addr_rom[  980] = 'h00000564; 	    d_addr_rom[  980] = 'h00000c38; 	    wdata_rom[  980] = 'h8b9c98ae; 	    wvalid_rom[  980] = 0; 
    i_addr_rom[  981] = 'h00000068; 	    d_addr_rom[  981] = 'h00000a70; 	    wdata_rom[  981] = 'hf3bad02d; 	    wvalid_rom[  981] = 1; 
    i_addr_rom[  982] = 'h0000026c; 	    d_addr_rom[  982] = 'h00000968; 	    wdata_rom[  982] = 'h79675dd5; 	    wvalid_rom[  982] = 1; 
    i_addr_rom[  983] = 'h0000069c; 	    d_addr_rom[  983] = 'h000008f8; 	    wdata_rom[  983] = 'h671a89de; 	    wvalid_rom[  983] = 1; 
    i_addr_rom[  984] = 'h00000518; 	    d_addr_rom[  984] = 'h00000c0c; 	    wdata_rom[  984] = 'h8fe16294; 	    wvalid_rom[  984] = 1; 
    i_addr_rom[  985] = 'h00000768; 	    d_addr_rom[  985] = 'h00000af4; 	    wdata_rom[  985] = 'hc193cf09; 	    wvalid_rom[  985] = 1; 
    i_addr_rom[  986] = 'h00000280; 	    d_addr_rom[  986] = 'h00000fe8; 	    wdata_rom[  986] = 'hb32c9c9a; 	    wvalid_rom[  986] = 0; 
    i_addr_rom[  987] = 'h0000075c; 	    d_addr_rom[  987] = 'h00000d34; 	    wdata_rom[  987] = 'h3dda23b8; 	    wvalid_rom[  987] = 1; 
    i_addr_rom[  988] = 'h0000038c; 	    d_addr_rom[  988] = 'h00000c4c; 	    wdata_rom[  988] = 'h33a5e677; 	    wvalid_rom[  988] = 1; 
    i_addr_rom[  989] = 'h00000730; 	    d_addr_rom[  989] = 'h0000088c; 	    wdata_rom[  989] = 'hdf88afaa; 	    wvalid_rom[  989] = 1; 
    i_addr_rom[  990] = 'h00000154; 	    d_addr_rom[  990] = 'h00000a80; 	    wdata_rom[  990] = 'hdf8921f2; 	    wvalid_rom[  990] = 0; 
    i_addr_rom[  991] = 'h000003e8; 	    d_addr_rom[  991] = 'h000008f8; 	    wdata_rom[  991] = 'hd22a54d8; 	    wvalid_rom[  991] = 0; 
    i_addr_rom[  992] = 'h000007dc; 	    d_addr_rom[  992] = 'h00000920; 	    wdata_rom[  992] = 'h23c0560b; 	    wvalid_rom[  992] = 0; 
    i_addr_rom[  993] = 'h00000614; 	    d_addr_rom[  993] = 'h00000f58; 	    wdata_rom[  993] = 'h64514c9f; 	    wvalid_rom[  993] = 1; 
    i_addr_rom[  994] = 'h000000dc; 	    d_addr_rom[  994] = 'h00000960; 	    wdata_rom[  994] = 'haa402afd; 	    wvalid_rom[  994] = 1; 
    i_addr_rom[  995] = 'h000007e4; 	    d_addr_rom[  995] = 'h0000094c; 	    wdata_rom[  995] = 'h07f8e524; 	    wvalid_rom[  995] = 0; 
    i_addr_rom[  996] = 'h00000310; 	    d_addr_rom[  996] = 'h00000904; 	    wdata_rom[  996] = 'h6f363563; 	    wvalid_rom[  996] = 0; 
    i_addr_rom[  997] = 'h000001a8; 	    d_addr_rom[  997] = 'h00000d74; 	    wdata_rom[  997] = 'h7cbc9026; 	    wvalid_rom[  997] = 1; 
    i_addr_rom[  998] = 'h00000738; 	    d_addr_rom[  998] = 'h00000a1c; 	    wdata_rom[  998] = 'ha1260194; 	    wvalid_rom[  998] = 0; 
    i_addr_rom[  999] = 'h00000660; 	    d_addr_rom[  999] = 'h00000fbc; 	    wdata_rom[  999] = 'hd5cf3ada; 	    wvalid_rom[  999] = 0; 
    i_addr_rom[ 1000] = 'h00000510; 	    d_addr_rom[ 1000] = 'h00000964; 	    wdata_rom[ 1000] = 'h8ceb6d18; 	    wvalid_rom[ 1000] = 1; 
    i_addr_rom[ 1001] = 'h00000628; 	    d_addr_rom[ 1001] = 'h00000ff0; 	    wdata_rom[ 1001] = 'hfd47d476; 	    wvalid_rom[ 1001] = 0; 
    i_addr_rom[ 1002] = 'h00000788; 	    d_addr_rom[ 1002] = 'h00000fdc; 	    wdata_rom[ 1002] = 'he87b542a; 	    wvalid_rom[ 1002] = 1; 
    i_addr_rom[ 1003] = 'h00000054; 	    d_addr_rom[ 1003] = 'h00000fa0; 	    wdata_rom[ 1003] = 'h831a995c; 	    wvalid_rom[ 1003] = 1; 
    i_addr_rom[ 1004] = 'h00000020; 	    d_addr_rom[ 1004] = 'h00000c38; 	    wdata_rom[ 1004] = 'h0b4f8f21; 	    wvalid_rom[ 1004] = 0; 
    i_addr_rom[ 1005] = 'h00000274; 	    d_addr_rom[ 1005] = 'h00000ee4; 	    wdata_rom[ 1005] = 'h0354ce45; 	    wvalid_rom[ 1005] = 0; 
    i_addr_rom[ 1006] = 'h0000003c; 	    d_addr_rom[ 1006] = 'h00000d0c; 	    wdata_rom[ 1006] = 'hc3f73ad7; 	    wvalid_rom[ 1006] = 1; 
    i_addr_rom[ 1007] = 'h0000031c; 	    d_addr_rom[ 1007] = 'h00000864; 	    wdata_rom[ 1007] = 'h9bf6a07c; 	    wvalid_rom[ 1007] = 1; 
    i_addr_rom[ 1008] = 'h000003d4; 	    d_addr_rom[ 1008] = 'h00000b20; 	    wdata_rom[ 1008] = 'hfd5c21ee; 	    wvalid_rom[ 1008] = 1; 
    i_addr_rom[ 1009] = 'h0000072c; 	    d_addr_rom[ 1009] = 'h00000aa0; 	    wdata_rom[ 1009] = 'hacdccfbf; 	    wvalid_rom[ 1009] = 0; 
    i_addr_rom[ 1010] = 'h0000070c; 	    d_addr_rom[ 1010] = 'h00000870; 	    wdata_rom[ 1010] = 'h5f0a9cad; 	    wvalid_rom[ 1010] = 0; 
    i_addr_rom[ 1011] = 'h000003a4; 	    d_addr_rom[ 1011] = 'h00000e2c; 	    wdata_rom[ 1011] = 'h0d35ea7f; 	    wvalid_rom[ 1011] = 0; 
    i_addr_rom[ 1012] = 'h000004b4; 	    d_addr_rom[ 1012] = 'h00000d68; 	    wdata_rom[ 1012] = 'hc8c00121; 	    wvalid_rom[ 1012] = 0; 
    i_addr_rom[ 1013] = 'h000001e0; 	    d_addr_rom[ 1013] = 'h00000f14; 	    wdata_rom[ 1013] = 'h31dbb89c; 	    wvalid_rom[ 1013] = 0; 
    i_addr_rom[ 1014] = 'h00000624; 	    d_addr_rom[ 1014] = 'h00000dc0; 	    wdata_rom[ 1014] = 'h818e5151; 	    wvalid_rom[ 1014] = 1; 
    i_addr_rom[ 1015] = 'h00000388; 	    d_addr_rom[ 1015] = 'h00000ca8; 	    wdata_rom[ 1015] = 'hcfef5b13; 	    wvalid_rom[ 1015] = 1; 
    i_addr_rom[ 1016] = 'h00000784; 	    d_addr_rom[ 1016] = 'h00000db4; 	    wdata_rom[ 1016] = 'h355cd9f9; 	    wvalid_rom[ 1016] = 0; 
    i_addr_rom[ 1017] = 'h00000234; 	    d_addr_rom[ 1017] = 'h00000e0c; 	    wdata_rom[ 1017] = 'hcba80e3b; 	    wvalid_rom[ 1017] = 0; 
    i_addr_rom[ 1018] = 'h000000ac; 	    d_addr_rom[ 1018] = 'h00000e78; 	    wdata_rom[ 1018] = 'h98eae9fb; 	    wvalid_rom[ 1018] = 0; 
    i_addr_rom[ 1019] = 'h00000494; 	    d_addr_rom[ 1019] = 'h00000b74; 	    wdata_rom[ 1019] = 'h44457704; 	    wvalid_rom[ 1019] = 0; 
    i_addr_rom[ 1020] = 'h000007cc; 	    d_addr_rom[ 1020] = 'h00000c20; 	    wdata_rom[ 1020] = 'he7743182; 	    wvalid_rom[ 1020] = 0; 
    i_addr_rom[ 1021] = 'h000000f8; 	    d_addr_rom[ 1021] = 'h00000ebc; 	    wdata_rom[ 1021] = 'h5e9baa30; 	    wvalid_rom[ 1021] = 0; 
    i_addr_rom[ 1022] = 'h000005b8; 	    d_addr_rom[ 1022] = 'h00000bb4; 	    wdata_rom[ 1022] = 'h29b82b9e; 	    wvalid_rom[ 1022] = 0; 
    i_addr_rom[ 1023] = 'h00000308; 	    d_addr_rom[ 1023] = 'h00000800; 	    wdata_rom[ 1023] = 'he4067be5; 	    wvalid_rom[ 1023] = 0; 

end
// for icache 
wire            i_rvalid_pipe;
wire            i_rready_pipe;
wire    [31:0]  i_raddr_pipe;
wire    [31:0]  i_rdata_pipe;
wire            i_rvalid;
wire            i_rready;
// icache && arbiter 
wire    [31:0]  i_raddr;
wire    [31:0]  i_rdata;
wire            i_rlast;
wire    [2:0]   i_rsize;
wire    [7:0]   i_rlen;
// icache_debug
reg             i_rvalid_ff;
reg     [31:0]  i_raddr_ff;
reg             i_error_reg;
reg             i_pass_reg;
wire    [31:0]  i_correct_data;

// for dcache
wire    [31:0]  d_addr_pipe;
wire            d_rvalid_pipe;
wire            d_rready_pipe;
wire    [31:0]  d_rdata_pipe;
wire            d_wvalid_pipe;
wire            d_wready_pipe;
wire    [31:0]  d_wdata_pipe;
wire    [3:0]   d_wstrb_pipe;
// dcache && arbiter
wire            d_rvalid;
wire            d_rready;
wire    [31:0]  d_raddr;
wire    [31:0]  d_rdata;
wire            d_rlast;
wire    [2:0]   d_rsize;
wire    [7:0]   d_rlen;
wire            d_wvalid;
wire            d_wready;
wire    [31:0]  d_waddr;
wire    [31:0]  d_wdata;
wire    [3:0]   d_wstrb;
wire            d_wlast;
wire    [2:0]   d_wsize;
wire    [7:0]   d_wlen;
wire            d_bvalid;
wire            d_bready;
// dcache_debug
reg             d_rvalid_ff;
reg             d_wvalid_ff;
reg     [31:0]  d_wdata_ff;
reg     [31:0]  d_addr_ff;
reg             d_error_reg;
reg             d_pass_reg;
wire    [31:0]  d_correct_data;

// arbiter with main mem
wire    [31:0]  araddr;
wire            arvalid;
wire            arready;
wire    [7:0]   arlen;
wire    [2:0]   arsize;
wire    [1:0]   arburst;
wire    [31:0]  rdata;
wire    [1:0]   rresp;
wire            rvalid;
wire            rready;
wire            rlast;
wire    [31:0]  awaddr;
wire            awvalid;
wire            awready;
wire    [7:0]   awlen;
wire    [2:0]   awsize;
wire    [1:0]   awburst;
wire    [31:0]  wdata;
wire    [3:0]   wstrb;
wire            wvalid;
wire            wready;
wire            wlast;
wire    [1:0]   bresp;
wire            bvalid;
wire            bready;

assign i_raddr_pipe = i_addr_rom[i_test_index];
assign i_correct_data = data_ram[i_raddr_ff >> 2];
assign i_rvalid_pipe = 1'b1;
// simulate IF1-IF2 register i_rvalid_ff && i_raddr_ff
always @(posedge clk) begin
    if(!rstn) begin
        i_rvalid_ff <= 0;
        i_raddr_ff <= 0;
    end
    else if(!(i_rvalid_ff && !i_rready_pipe))begin
        i_rvalid_ff <= i_rvalid_pipe;
        i_raddr_ff <= i_raddr_pipe;
    end
end
// update i_test_index
always @(posedge clk) begin
    if(!rstn) begin
        i_test_index <= 0;
        i_pass_reg <= 0;
    end
    else if (i_test_index >= (TOTAL_WORD_NUM / 2-1)) begin
        i_test_index <= (TOTAL_WORD_NUM / 2-1);
        i_pass_reg <= 1;
    end
    else if(!(i_rvalid_ff && !i_rready_pipe) && !i_error_reg) begin
        i_test_index <= i_test_index + 1;
    end
end
// update i_error 
always @(posedge clk) begin
    if(!rstn) begin
        i_error_reg <= 0;
    end
    else if(i_error_reg) begin
        i_error_reg <= 1;
    end
    else if(i_rvalid_ff && i_rready_pipe) begin
        i_error_reg <= !(i_rdata_pipe  == i_correct_data);
    end
end

assign d_addr_pipe           = d_addr_rom[d_test_index];
assign d_correct_data   = data_ram[d_addr_ff >> 2];
assign d_rvalid_pipe         = !wvalid_rom[d_test_index];
assign d_wvalid_pipe         = wvalid_rom[d_test_index];
assign d_wdata_pipe          = wdata_rom[d_test_index];
assign d_wstrb_pipe          = d_wvalid_pipe ? 4'b1111 : 4'b0000;
// simulate EX-MEM register
always @(posedge clk) begin
    if(!rstn) begin
        d_rvalid_ff <= 0;
        d_addr_ff   <= 0;
        d_wvalid_ff <= 0;
        d_wdata_ff  <= 0;
    end
    else if(!(d_rvalid_ff && !d_rready_pipe) && !(d_wvalid_ff && !d_wready_pipe))begin
        d_rvalid_ff <= d_rvalid_pipe;
        d_addr_ff   <= d_addr_pipe;
        d_wvalid_ff <= d_wvalid_pipe;
        d_wdata_ff  <= d_wdata_pipe;
    end
end
// update d_test_index
always @(posedge clk) begin
    if(!rstn) begin
        d_test_index    <= TOTAL_WORD_NUM / 2;
        d_pass_reg      <= 0;
    end
    else if (d_test_index >= (TOTAL_WORD_NUM-1)) begin
        d_test_index    <= (TOTAL_WORD_NUM-1);
        d_pass_reg      <= 1;
    end
    else if(!(d_rvalid_ff && !d_rready_pipe)  && !(d_wvalid_ff && !d_wready_pipe) && !d_error_reg) begin
        d_test_index    <= d_test_index + 1;
    end
end
// update data_ram
always @(posedge clk) begin
    if(d_wvalid_ff && d_wready_pipe) begin
        data_ram[d_addr_ff >> 2] <= d_wdata_ff;
    end
end
// update d_error 
always @(posedge clk) begin
    if(!rstn) begin
        d_error_reg <= 0;
    end
    else if(d_error_reg) begin
        d_error_reg <= 1;
    end
    else if(d_rvalid_ff && d_rready_pipe) begin
        d_error_reg <= !(d_rdata_pipe  == d_correct_data);
    end
end

icache #(
  .INDEX_WIDTH          (INDEX_WIDTH),
  .WORD_OFFSET_WIDTH    (WORD_OFFSET_WIDTH)
)
icache_dut (
    .clk      (clk ),
    .rstn     (rstn ),
    .rvalid   (i_rvalid_pipe ),
    .rready   (i_rready_pipe ),
    .raddr    (i_raddr_pipe ),
    .rdata    (i_rdata_pipe ),

    .i_rvalid (i_rvalid ),
    .i_rready (i_rready ),
    .i_raddr  (i_raddr ),
    .i_rdata  (i_rdata ),
    .i_rlast  (i_rlast ),
    .i_rsize  (i_rsize ),
    .i_rlen   (i_rlen)
);
dcache #(
    .INDEX_WIDTH        (INDEX_WIDTH ),
    .WORD_OFFSET_WIDTH  (WORD_OFFSET_WIDTH )
)
dcache_dut (
    .clk      (clk ),
    .rstn     (rstn ),
    .addr     (d_addr_pipe ),
    .rvalid   (d_rvalid_pipe ),
    .rready   (d_rready_pipe ),
    .rdata    (d_rdata_pipe ),
    .wvalid   (d_wvalid_pipe ),
    .wready   (d_wready_pipe ),
    .wdata    (d_wdata_pipe ),
    .wstrb    (d_wstrb_pipe ),
    .d_rvalid (d_rvalid ),
    .d_rready (d_rready ),
    .d_raddr  (d_raddr ),
    .d_rdata  (d_rdata ),
    .d_rlast  (d_rlast ),
    .d_rsize  (d_rsize ),
    .d_rlen   (d_rlen ),
    .d_wvalid (d_wvalid ),
    .d_wready (d_wready ),
    .d_waddr  (d_waddr ),
    .d_wdata  (d_wdata ),
    .d_wstrb  (d_wstrb ),
    .d_wlast  (d_wlast ),
    .d_wsize  (d_wsize ),
    .d_wlen   (d_wlen ),
    .d_bvalid (d_bvalid ),
    .d_bready (d_bready )
);

axi_arbiter axi_arbiter_dut (
    .clk      (clk ),
    .rstn     (rstn ),
    .i_rvalid (i_rvalid ),
    .i_rready (i_rready ),
    .i_raddr  (i_raddr ),
    .i_rdata  (i_rdata ),
    .i_rlast  (i_rlast ),
    .i_rsize  (i_rsize ),
    .i_rlen   (i_rlen ),
    .d_rvalid (d_rvalid ),
    .d_rready (d_rready ),
    .d_raddr  (d_raddr ),
    .d_rdata  (d_rdata ),
    .d_rlast  (d_rlast ),
    .d_rsize  (d_rsize ),
    .d_rlen   (d_rlen ),
    .d_wvalid (d_wvalid ),
    .d_wready (d_wready ),
    .d_waddr  (d_waddr ),
    .d_wdata  (d_wdata ),
    .d_wstrb  (d_wstrb ),
    .d_wlast  (d_wlast ),
    .d_wsize  (d_wsize ),
    .d_wlen   (d_wlen ),
    .d_bvalid (d_bvalid ),
    .d_bready (d_bready ),
    .araddr   (araddr ),
    .arvalid  (arvalid ),
    .arready  (arready ),
    .arlen    (arlen ),
    .arsize   (arsize ),
    .arburst  (arburst ),
    .rdata    (rdata ),
    .rresp    (rresp ),
    .rvalid   (rvalid ),
    .rready   (rready ),
    .rlast    (rlast ),
    .awaddr   (awaddr ),
    .awvalid  (awvalid ),
    .awready  (awready ),
    .awlen    (awlen ),
    .awsize   (awsize ),
    .awburst  (awburst ),
    .wdata    (wdata ),
    .wstrb    (wstrb ),
    .wvalid   (wvalid ),
    .wready   (wready ),
    .wlast    (wlast ),
    .bresp    (bresp ),
    .bvalid   (bvalid ),
    .bready   (bready)
);
main_memory main_mem(
    .s_aclk         (clk ),
    .s_aresetn      (rstn ),
    .s_axi_araddr   (araddr ),
    .s_axi_arburst  (arburst ),
    .s_axi_arid     (4'b0),
    .s_axi_arlen    (arlen ),
    .s_axi_arready  (arready ),
    .s_axi_arsize   (arsize ),
    .s_axi_arvalid  (arvalid ),
    .s_axi_awaddr   (awaddr ),
    .s_axi_awburst  (awburst ),
    .s_axi_awid     (4'b0),
    .s_axi_awlen    (awlen ),
    .s_axi_awready  (awready ),
    .s_axi_awsize   (awsize ),
    .s_axi_awvalid  (awvalid ),
    .s_axi_bid      (),
    .s_axi_bready   (bready ),
    .s_axi_bresp    (bresp ),
    .s_axi_bvalid   (bvalid ),
    .s_axi_rdata    (rdata ),
    .s_axi_rid      (),
    .s_axi_rlast    (rlast ),
    .s_axi_rready   (rready ),
    .s_axi_rresp    (rresp ),
    .s_axi_rvalid   (rvalid ),
    .s_axi_wdata    (wdata ),
    .s_axi_wlast    (wlast ),
    .s_axi_wready   (wready ),
    .s_axi_wstrb    (wstrb ),
    .s_axi_wvalid   (wvalid )
);
endmodule

